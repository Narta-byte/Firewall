library IEEE;
library std;
use IEEE.std_logic_1164.all;
use IEEE.NUMERIC_STD.all;

entity input_packet_rom is
  port (
    address : in std_logic_vector(12 downto 0);
    data_out : out std_logic_vector(9 downto 0) 
  );
end entity;


architecture input_packet_rom_arch of input_packet_rom is
    type ROM_type is array (0 to 5599) of std_logic_vector(9 downto 0);

    constant ROM : ROM_type := (0 => "1001110000",
                                1 => "1011011000",
                                2 => "1101000000",
                                3 => "0001011100",
                                4 => "0100101100",
                                5 => "0000100100",
                                6 => "0110000000",
                                7 => "0011001000",
                                8 => "1011000100",
                                9 => "1000110000",
                                10 => "0100011100",
                                11 => "0100111100",
                                12 => "0000100000",
                                13 => "0000000000",
                                14 => "0100010101",
                                15 => "0100010110",
                                16 => "0000000000",
                                17 => "0000000000",
                                18 => "0011000000",
                                19 => "0000000000",
                                20 => "0000000000",
                                21 => "0100000000",
                                22 => "0000000000",
                                23 => "0011000100",
                                24 => "0000011000",
                                25 => "0111110100",
                                26 => "1001101000",
                                27 => "1011100100",
                                28 => "1001111100",
                                29 => "0101000000",
                                30 => "1000000000",
                                31 => "1100000000",
                                32 => "1010100000",
                                33 => "0000000100",
                                34 => "0110011000",
                                35 => "0001111100",
                                36 => "1001110000",
                                37 => "1110010000",
                                38 => "1100010000",
                                39 => "0100110000",
                                40 => "0010000000",
                                41 => "0101101000",
                                42 => "1010101000",
                                43 => "0110011000",
                                44 => "1001001100",
                                45 => "0111110100",
                                46 => "0110110100",
                                47 => "0111000000",
                                48 => "0001001000",
                                49 => "1010010100",
                                50 => "0110010000",
                                51 => "1000001000",
                                52 => "0101000000",
                                53 => "0000000000",
                                54 => "0000000000",
                                55 => "0000001000",
                                56 => "0000010000",
                                57 => "0000010100",
                                58 => "1011010000",
                                59 => "0000000100",
                                60 => "0000000100",
                                61 => "0000010000",
                                62 => "0000001000",
                                63 => "1001110000",
                                64 => "1011011000",
                                65 => "1101000000",
                                66 => "0001011100",
                                67 => "0100101100",
                                68 => "0000100100",
                                69 => "0110000000",
                                70 => "0011001000",
                                71 => "1011000100",
                                72 => "1000110000",
                                73 => "0100011100",
                                74 => "0100111100",
                                75 => "0000100000",
                                76 => "0000000000",
                                77 => "0100010101",
                                78 => "0100010110",
                                79 => "0000000000",
                                80 => "0000000000",
                                81 => "0011000000",
                                82 => "0000000000",
                                83 => "0000000000",
                                84 => "0100000000",
                                85 => "0000000000",
                                86 => "0011001000",
                                87 => "0000011000",
                                88 => "1011100100",
                                89 => "0000010100",
                                90 => "0101111000",
                                91 => "1110110100",
                                92 => "0110111000",
                                93 => "1100011100",
                                94 => "1100000000",
                                95 => "1010100000",
                                96 => "0000000100",
                                97 => "0110011000",
                                98 => "0000000100",
                                99 => "1011101100",
                                100 => "1110010000",
                                101 => "1100010100",
                                102 => "1011111100",
                                103 => "0111111000",
                                104 => "0100010100",
                                105 => "1001010000",
                                106 => "1111101100",
                                107 => "0001010000",
                                108 => "1101101000",
                                109 => "0111010100",
                                110 => "0111000000",
                                111 => "0001001000",
                                112 => "1111101000",
                                113 => "1111000000",
                                114 => "0011011100",
                                115 => "0011110100",
                                116 => "0000000000",
                                117 => "0000000000",
                                118 => "0000001000",
                                119 => "0000010000",
                                120 => "0000010100",
                                121 => "1011010000",
                                122 => "0000000100",
                                123 => "0000000100",
                                124 => "0000010000",
                                125 => "0000001000",
                                126 => "1001110000",
                                127 => "1011011000",
                                128 => "1101000000",
                                129 => "0001011100",
                                130 => "0100101100",
                                131 => "0000100100",
                                132 => "0110000000",
                                133 => "0011001000",
                                134 => "1011000100",
                                135 => "1000110000",
                                136 => "0100011100",
                                137 => "0100111100",
                                138 => "0000100000",
                                139 => "0000000000",
                                140 => "0100010101",
                                141 => "0100010110",
                                142 => "0000000000",
                                143 => "0000000000",
                                144 => "0011000000",
                                145 => "0000000000",
                                146 => "0000000000",
                                147 => "0100000000",
                                148 => "0000000000",
                                149 => "0011001000",
                                150 => "0000011000",
                                151 => "1011100100",
                                152 => "0000010100",
                                153 => "0101111000",
                                154 => "1110110100",
                                155 => "0110111000",
                                156 => "1100011100",
                                157 => "1100000000",
                                158 => "1010100000",
                                159 => "0000000100",
                                160 => "0110011000",
                                161 => "0000000100",
                                162 => "1011101100",
                                163 => "1110010000",
                                164 => "1100011000",
                                165 => "1110110100",
                                166 => "1111011100",
                                167 => "0010110000",
                                168 => "1001011000",
                                169 => "1010011100",
                                170 => "1011001100",
                                171 => "0100011100",
                                172 => "1111110000",
                                173 => "0111000000",
                                174 => "0001001000",
                                175 => "1111101000",
                                176 => "1111000000",
                                177 => "0000011100",
                                178 => "1001110000",
                                179 => "0000000000",
                                180 => "0000000000",
                                181 => "0000001000",
                                182 => "0000010000",
                                183 => "0000010100",
                                184 => "1011010000",
                                185 => "0000000100",
                                186 => "0000000100",
                                187 => "0000010000",
                                188 => "0000001000",
                                189 => "1001110000",
                                190 => "1011011000",
                                191 => "1101000000",
                                192 => "0001011100",
                                193 => "0100101100",
                                194 => "0000100100",
                                195 => "0110000000",
                                196 => "0011001000",
                                197 => "1011000100",
                                198 => "1000110000",
                                199 => "0100011100",
                                200 => "0100111100",
                                201 => "0000100000",
                                202 => "0000000000",
                                203 => "0100010101",
                                204 => "0100010110",
                                205 => "0000000000",
                                206 => "0000000000",
                                207 => "0011000000",
                                208 => "1110111000",
                                209 => "1110100100",
                                210 => "0100000000",
                                211 => "0000000000",
                                212 => "0111011000",
                                213 => "0000011000",
                                214 => "0101000000",
                                215 => "0011100000",
                                216 => "0000110100",
                                217 => "0110101100",
                                218 => "1111011000",
                                219 => "0010110000",
                                220 => "1100000000",
                                221 => "1010100000",
                                222 => "0000000100",
                                223 => "0110011000",
                                224 => "0000000100",
                                225 => "1011101100",
                                226 => "1110010000",
                                227 => "1100011100",
                                228 => "0011101100",
                                229 => "0111101100",
                                230 => "1001100000",
                                231 => "1110111000",
                                232 => "1111010100",
                                233 => "0110110100",
                                234 => "0011001100",
                                235 => "0010011000",
                                236 => "0111000000",
                                237 => "0001001000",
                                238 => "1111101000",
                                239 => "1111000000",
                                240 => "1101111100",
                                241 => "0000101100",
                                242 => "0000000000",
                                243 => "0000000000",
                                244 => "0000001000",
                                245 => "0000010000",
                                246 => "0000010100",
                                247 => "1010000000",
                                248 => "0000000100",
                                249 => "0000000100",
                                250 => "0000010000",
                                251 => "0000001000",
                                252 => "1001110000",
                                253 => "1011011000",
                                254 => "1101000000",
                                255 => "0001011100",
                                256 => "0100101100",
                                257 => "0000100100",
                                258 => "0110000000",
                                259 => "0011001000",
                                260 => "1011000100",
                                261 => "1000110000",
                                262 => "0100011100",
                                263 => "0100111100",
                                264 => "0000100000",
                                265 => "0000000000",
                                266 => "0100010101",
                                267 => "0100010110",
                                268 => "0000000000",
                                269 => "0000000000",
                                270 => "0011000000",
                                271 => "0000000000",
                                272 => "0000000000",
                                273 => "0100000000",
                                274 => "0000000000",
                                275 => "0011000100",
                                276 => "0000011000",
                                277 => "0111110100",
                                278 => "1001101000",
                                279 => "1011100100",
                                280 => "1001111100",
                                281 => "0101000000",
                                282 => "1000000000",
                                283 => "1100000000",
                                284 => "1010100000",
                                285 => "0000000100",
                                286 => "0110011000",
                                287 => "0001111100",
                                288 => "1001110000",
                                289 => "1110010000",
                                290 => "1100100000",
                                291 => "1010100000",
                                292 => "0000010000",
                                293 => "1001111100",
                                294 => "0111111100",
                                295 => "1001101000",
                                296 => "0011000000",
                                297 => "1100100000",
                                298 => "0010111100",
                                299 => "0111000000",
                                300 => "0001001000",
                                301 => "1010010100",
                                302 => "0110010000",
                                303 => "0110001100",
                                304 => "0011001100",
                                305 => "0000000000",
                                306 => "0000000000",
                                307 => "0000001000",
                                308 => "0000010000",
                                309 => "0000010100",
                                310 => "1011010000",
                                311 => "0000000100",
                                312 => "0000000100",
                                313 => "0000010000",
                                314 => "0000001000",
                                315 => "1001110000",
                                316 => "1011011000",
                                317 => "1101000000",
                                318 => "0001011100",
                                319 => "0100101100",
                                320 => "0000100100",
                                321 => "0110000000",
                                322 => "0011001000",
                                323 => "1011000100",
                                324 => "1000110000",
                                325 => "0100011100",
                                326 => "0100111100",
                                327 => "0000100000",
                                328 => "0000000000",
                                329 => "0100010101",
                                330 => "0100010110",
                                331 => "0000000000",
                                332 => "0000000000",
                                333 => "0011000000",
                                334 => "0000000000",
                                335 => "0000000000",
                                336 => "0100000000",
                                337 => "0000000000",
                                338 => "0011001000",
                                339 => "0000011000",
                                340 => "0111110000",
                                341 => "0011001100",
                                342 => "0101101100",
                                343 => "1100011000",
                                344 => "1010111000",
                                345 => "1100000000",
                                346 => "1100000000",
                                347 => "1010100000",
                                348 => "0000000100",
                                349 => "0110011000",
                                350 => "0000000100",
                                351 => "1011101100",
                                352 => "1110010000",
                                353 => "1100100100",
                                354 => "1100111100",
                                355 => "0111100100",
                                356 => "0110000000",
                                357 => "0010001000",
                                358 => "1001010000",
                                359 => "0010101000",
                                360 => "1011100000",
                                361 => "1111000100",
                                362 => "0111000000",
                                363 => "0001001000",
                                364 => "1010010100",
                                365 => "0110010000",
                                366 => "1010110100",
                                367 => "1111000000",
                                368 => "0000000000",
                                369 => "0000000000",
                                370 => "0000001000",
                                371 => "0000010000",
                                372 => "0000010100",
                                373 => "1001110000",
                                374 => "0000000100",
                                375 => "0000000100",
                                376 => "0000010000",
                                377 => "0000001000",
                                378 => "1001110000",
                                379 => "1011011000",
                                380 => "1101000000",
                                381 => "0001011100",
                                382 => "0100101100",
                                383 => "0000100100",
                                384 => "0110000000",
                                385 => "0011001000",
                                386 => "1011000100",
                                387 => "1000110000",
                                388 => "0100011100",
                                389 => "0100111100",
                                390 => "0000100000",
                                391 => "0000000000",
                                392 => "0100010101",
                                393 => "0100010110",
                                394 => "0000000000",
                                395 => "0000000000",
                                396 => "0011000000",
                                397 => "0000000000",
                                398 => "0000000000",
                                399 => "0100000000",
                                400 => "0000000000",
                                401 => "0011001000",
                                402 => "0000011000",
                                403 => "0111110000",
                                404 => "0010001100",
                                405 => "0101101100",
                                406 => "1100011000",
                                407 => "1010111000",
                                408 => "1101000000",
                                409 => "1100000000",
                                410 => "1010100000",
                                411 => "0000000100",
                                412 => "0110011000",
                                413 => "0000000100",
                                414 => "1011101100",
                                415 => "1110010000",
                                416 => "1100101000",
                                417 => "0111101000",
                                418 => "0000011100",
                                419 => "0101011000",
                                420 => "0100010100",
                                421 => "1111111000",
                                422 => "1101101000",
                                423 => "0010000000",
                                424 => "0100100100",
                                425 => "0111000000",
                                426 => "0001001000",
                                427 => "1010010100",
                                428 => "0110010000",
                                429 => "0011101100",
                                430 => "0010011100",
                                431 => "0000000000",
                                432 => "0000000000",
                                433 => "0000001000",
                                434 => "0000010000",
                                435 => "0000010100",
                                436 => "1001110000",
                                437 => "0000000100",
                                438 => "0000000100",
                                439 => "0000010000",
                                440 => "0000001000",
                                441 => "1001110000",
                                442 => "1011011000",
                                443 => "1101000000",
                                444 => "0001011100",
                                445 => "0100101100",
                                446 => "0000100100",
                                447 => "0110000000",
                                448 => "0011001000",
                                449 => "1011000100",
                                450 => "1000110000",
                                451 => "0100011100",
                                452 => "0100111100",
                                453 => "0000100000",
                                454 => "0000000000",
                                455 => "0100010101",
                                456 => "0100010110",
                                457 => "0000000000",
                                458 => "0000000000",
                                459 => "0011000000",
                                460 => "0000000000",
                                461 => "0000000000",
                                462 => "0100000000",
                                463 => "0000000000",
                                464 => "0011000100",
                                465 => "0000011000",
                                466 => "0111110100",
                                467 => "1001101000",
                                468 => "1011100100",
                                469 => "1001111100",
                                470 => "0101000000",
                                471 => "1000000000",
                                472 => "1100000000",
                                473 => "1010100000",
                                474 => "0000000100",
                                475 => "0110011000",
                                476 => "0001111100",
                                477 => "1001110000",
                                478 => "1110010000",
                                479 => "1100101100",
                                480 => "1000110100",
                                481 => "0011000000",
                                482 => "0110001000",
                                483 => "0111001100",
                                484 => "0111111000",
                                485 => "0000101100",
                                486 => "0101101100",
                                487 => "1111100000",
                                488 => "0111000000",
                                489 => "0001001000",
                                490 => "1010010100",
                                491 => "0110010000",
                                492 => "0100001100",
                                493 => "0110110100",
                                494 => "0000000000",
                                495 => "0000000000",
                                496 => "0000001000",
                                497 => "0000010000",
                                498 => "0000010100",
                                499 => "1011010000",
                                500 => "0000000100",
                                501 => "0000000100",
                                502 => "0000010000",
                                503 => "0000001000",
                                504 => "1001110000",
                                505 => "1011011000",
                                506 => "1101000000",
                                507 => "0001011100",
                                508 => "0100101100",
                                509 => "0000100100",
                                510 => "0110000000",
                                511 => "0011001000",
                                512 => "1011000100",
                                513 => "1000110000",
                                514 => "0100011100",
                                515 => "0100111100",
                                516 => "0000100000",
                                517 => "0000000000",
                                518 => "0100010101",
                                519 => "0100010110",
                                520 => "1000000000",
                                521 => "0000000000",
                                522 => "0011000000",
                                523 => "1101111000",
                                524 => "1000011100",
                                525 => "0000000000",
                                526 => "0000000000",
                                527 => "0111011000",
                                528 => "0000011000",
                                529 => "0000101100",
                                530 => "0001101000",
                                531 => "1000111000",
                                532 => "1111101100",
                                533 => "0000100100",
                                534 => "1001110100",
                                535 => "1100000000",
                                536 => "1010100000",
                                537 => "0000000100",
                                538 => "0110011000",
                                539 => "0000000100",
                                540 => "1011101100",
                                541 => "1110010000",
                                542 => "1100110100",
                                543 => "1101011000",
                                544 => "0001000100",
                                545 => "0010001100",
                                546 => "1011101000",
                                547 => "1111111000",
                                548 => "1101110100",
                                549 => "1000110100",
                                550 => "0001010100",
                                551 => "0111000000",
                                552 => "0001001000",
                                553 => "1111111100",
                                554 => "1111111100",
                                555 => "1011110000",
                                556 => "0011111000",
                                557 => "0000000000",
                                558 => "0000000000",
                                559 => "0000001000",
                                560 => "0000010000",
                                561 => "0000010100",
                                562 => "1001011000",
                                563 => "0000000100",
                                564 => "0000000100",
                                565 => "0000010000",
                                566 => "0000001000",
                                567 => "1001110000",
                                568 => "1011011000",
                                569 => "1101000000",
                                570 => "0001011100",
                                571 => "0100101100",
                                572 => "0000100100",
                                573 => "0110000000",
                                574 => "0011001000",
                                575 => "1011000100",
                                576 => "1000110000",
                                577 => "0100011100",
                                578 => "0100111100",
                                579 => "0000100000",
                                580 => "0000000000",
                                581 => "0100010101",
                                582 => "0100010110",
                                583 => "0000000000",
                                584 => "0000000000",
                                585 => "0011000000",
                                586 => "0000000000",
                                587 => "0000000000",
                                588 => "0100000000",
                                589 => "0000000000",
                                590 => "1101101000",
                                591 => "0000011000",
                                592 => "0101111000",
                                593 => "0111011000",
                                594 => "0001001000",
                                595 => "1101100000",
                                596 => "0110110100",
                                597 => "0110101100",
                                598 => "1100000000",
                                599 => "1010100000",
                                600 => "0000000100",
                                601 => "0110011000",
                                602 => "0000000100",
                                603 => "1011101100",
                                604 => "1110010000",
                                605 => "1100110000",
                                606 => "1110100000",
                                607 => "0100100000",
                                608 => "0000011100",
                                609 => "0111011100",
                                610 => "0010101000",
                                611 => "1010000100",
                                612 => "1101101100",
                                613 => "1010010100",
                                614 => "0111000000",
                                615 => "0001001000",
                                616 => "0110100100",
                                617 => "0000001100",
                                618 => "1111101100",
                                619 => "0010101100",
                                620 => "0000000000",
                                621 => "0000000000",
                                622 => "0000001000",
                                623 => "0000010000",
                                624 => "0000010100",
                                625 => "1011010000",
                                626 => "0000000100",
                                627 => "0000000100",
                                628 => "0000010000",
                                629 => "0000001000",
                                630 => "1001110000",
                                631 => "1011011000",
                                632 => "1101000000",
                                633 => "0001011100",
                                634 => "0100101100",
                                635 => "0000100100",
                                636 => "0110000000",
                                637 => "0011001000",
                                638 => "1011000100",
                                639 => "1000110000",
                                640 => "0100011100",
                                641 => "0100111100",
                                642 => "0000100000",
                                643 => "0000000000",
                                644 => "0100010101",
                                645 => "0100010110",
                                646 => "0000000000",
                                647 => "0000000000",
                                648 => "0011000000",
                                649 => "0000000000",
                                650 => "0000000000",
                                651 => "0100000000",
                                652 => "0000000000",
                                653 => "0011100100",
                                654 => "0000011000",
                                655 => "0101110100",
                                656 => "0110111000",
                                657 => "0110100000",
                                658 => "0001001000",
                                659 => "1011101000",
                                660 => "0011100100",
                                661 => "1100000000",
                                662 => "1010100000",
                                663 => "0000000100",
                                664 => "0110011000",
                                665 => "0000000100",
                                666 => "1011101100",
                                667 => "1110010000",
                                668 => "1100111000",
                                669 => "1101011000",
                                670 => "1101001100",
                                671 => "0101111000",
                                672 => "1001011100",
                                673 => "0100110100",
                                674 => "0110101100",
                                675 => "0111100000",
                                676 => "1011001000",
                                677 => "0111000000",
                                678 => "0001001000",
                                679 => "1111111100",
                                680 => "1111111100",
                                681 => "1011110000",
                                682 => "1101111000",
                                683 => "0000000000",
                                684 => "0000000000",
                                685 => "0000001000",
                                686 => "0000010000",
                                687 => "0000010100",
                                688 => "0111100000",
                                689 => "0000000100",
                                690 => "0000000100",
                                691 => "0000010000",
                                692 => "0000001000",
                                693 => "1001110000",
                                694 => "1011011000",
                                695 => "1101000000",
                                696 => "0001011100",
                                697 => "0100101100",
                                698 => "0000100100",
                                699 => "0110000000",
                                700 => "0011001000",
                                701 => "1011000100",
                                702 => "1000110000",
                                703 => "0100011100",
                                704 => "0100111100",
                                705 => "0000100000",
                                706 => "0000000000",
                                707 => "0100010101",
                                708 => "0100010110",
                                709 => "0000000000",
                                710 => "0000000000",
                                711 => "0011000000",
                                712 => "0000000000",
                                713 => "0000000000",
                                714 => "0100000000",
                                715 => "0000000000",
                                716 => "0011000100",
                                717 => "0000011000",
                                718 => "0111110100",
                                719 => "1001101000",
                                720 => "1011100100",
                                721 => "1001111100",
                                722 => "0101000000",
                                723 => "1000000000",
                                724 => "1100000000",
                                725 => "1010100000",
                                726 => "0000000100",
                                727 => "0110011000",
                                728 => "0001111100",
                                729 => "1001110000",
                                730 => "1110010000",
                                731 => "1100111100",
                                732 => "1110011000",
                                733 => "0000101100",
                                734 => "1111011000",
                                735 => "0011100000",
                                736 => "1100100000",
                                737 => "0100010000",
                                738 => "1111110100",
                                739 => "1111110000",
                                740 => "0111000000",
                                741 => "0001001000",
                                742 => "1010010100",
                                743 => "0110010000",
                                744 => "0110101000",
                                745 => "1000101000",
                                746 => "0000000000",
                                747 => "0000000000",
                                748 => "0000001000",
                                749 => "0000010000",
                                750 => "0000010100",
                                751 => "1011010000",
                                752 => "0000000100",
                                753 => "0000000100",
                                754 => "0000010000",
                                755 => "0000001000",
                                756 => "1001110000",
                                757 => "1011011000",
                                758 => "1101000000",
                                759 => "0001011100",
                                760 => "0100101100",
                                761 => "0000100100",
                                762 => "0110000000",
                                763 => "0011001000",
                                764 => "1011000100",
                                765 => "1000110000",
                                766 => "0100011100",
                                767 => "0100111100",
                                768 => "0000100000",
                                769 => "0000000000",
                                770 => "0100010101",
                                771 => "0100010110",
                                772 => "0000000000",
                                773 => "0000000000",
                                774 => "0011000000",
                                775 => "0010001100",
                                776 => "1001000100",
                                777 => "0000000000",
                                778 => "0000000000",
                                779 => "1111010000",
                                780 => "0000011000",
                                781 => "0101110000",
                                782 => "1110001000",
                                783 => "1000111100",
                                784 => "1100110000",
                                785 => "1111010000",
                                786 => "0111100100",
                                787 => "1100000000",
                                788 => "1010100000",
                                789 => "0000000100",
                                790 => "0110011000",
                                791 => "0000000100",
                                792 => "1011101100",
                                793 => "1110010000",
                                794 => "1101001100",
                                795 => "0000101100",
                                796 => "0101100000",
                                797 => "1110101100",
                                798 => "1100000000",
                                799 => "0100001100",
                                800 => "0100110100",
                                801 => "0011000000",
                                802 => "1010100000",
                                803 => "0111000000",
                                804 => "0001001000",
                                805 => "0000010100",
                                806 => "1010000000",
                                807 => "1110010100",
                                808 => "1001000100",
                                809 => "0000000000",
                                810 => "0000000000",
                                811 => "0000001000",
                                812 => "0000010000",
                                813 => "0000010100",
                                814 => "1010000000",
                                815 => "0000000100",
                                816 => "0000000100",
                                817 => "0000010000",
                                818 => "0000001000",
                                819 => "1001110000",
                                820 => "1011011000",
                                821 => "1101000000",
                                822 => "0001011100",
                                823 => "0100101100",
                                824 => "0000100100",
                                825 => "0110000000",
                                826 => "0011001000",
                                827 => "1011000100",
                                828 => "1000110000",
                                829 => "0100011100",
                                830 => "0100111100",
                                831 => "0000100000",
                                832 => "0000000000",
                                833 => "0100010101",
                                834 => "0100010110",
                                835 => "0000000000",
                                836 => "0000000000",
                                837 => "0011000000",
                                838 => "0000000000",
                                839 => "0000000000",
                                840 => "0100000000",
                                841 => "0000000000",
                                842 => "0011100000",
                                843 => "0000011000",
                                844 => "1000110000",
                                845 => "1001111100",
                                846 => "0100010100",
                                847 => "0001000000",
                                848 => "1010111100",
                                849 => "0000101000",
                                850 => "1100000000",
                                851 => "1010100000",
                                852 => "0000000100",
                                853 => "0110011000",
                                854 => "0000000100",
                                855 => "1011101100",
                                856 => "1110010000",
                                857 => "1101001000",
                                858 => "1010110000",
                                859 => "0001100000",
                                860 => "0101001100",
                                861 => "1001000000",
                                862 => "0000001000",
                                863 => "1110100100",
                                864 => "1101101000",
                                865 => "1010100000",
                                866 => "0111000000",
                                867 => "0001001000",
                                868 => "1111111100",
                                869 => "1111111100",
                                870 => "0000100100",
                                871 => "0001111000",
                                872 => "0000000000",
                                873 => "0000000000",
                                874 => "0000001000",
                                875 => "0000010000",
                                876 => "0000010100",
                                877 => "1011010000",
                                878 => "0000000100",
                                879 => "0000000100",
                                880 => "0000010000",
                                881 => "0000001000",
                                882 => "1001110000",
                                883 => "1011011000",
                                884 => "1101000000",
                                885 => "0001011100",
                                886 => "0100101100",
                                887 => "0000100100",
                                888 => "0110000000",
                                889 => "0011001000",
                                890 => "1011000100",
                                891 => "1000110000",
                                892 => "0100011100",
                                893 => "0100111100",
                                894 => "0000100000",
                                895 => "0000000000",
                                896 => "0100010101",
                                897 => "0100010110",
                                898 => "0000000000",
                                899 => "0000000000",
                                900 => "0011000000",
                                901 => "1001110100",
                                902 => "1101110100",
                                903 => "0000000000",
                                904 => "0000000000",
                                905 => "1111001100",
                                906 => "0000011000",
                                907 => "1110010000",
                                908 => "0000010000",
                                909 => "1000111100",
                                910 => "1100110000",
                                911 => "1111010000",
                                912 => "0000101000",
                                913 => "1100000000",
                                914 => "1010100000",
                                915 => "0000000100",
                                916 => "0110011000",
                                917 => "0000000100",
                                918 => "1011101100",
                                919 => "1110010000",
                                920 => "1101010000",
                                921 => "0110100000",
                                922 => "1101111100",
                                923 => "1111001000",
                                924 => "0010110000",
                                925 => "1101110100",
                                926 => "1111010100",
                                927 => "1001011100",
                                928 => "0001100100",
                                929 => "0111000000",
                                930 => "0001001000",
                                931 => "0000010100",
                                932 => "1010000000",
                                933 => "1000000000",
                                934 => "1111001000",
                                935 => "0000000000",
                                936 => "0000000000",
                                937 => "0000001000",
                                938 => "0000010000",
                                939 => "0000010100",
                                940 => "1010000000",
                                941 => "0000000100",
                                942 => "0000000100",
                                943 => "0000010000",
                                944 => "0000001000",
                                945 => "1001110000",
                                946 => "1011011000",
                                947 => "1101000000",
                                948 => "0001011100",
                                949 => "0100101100",
                                950 => "0000100100",
                                951 => "0110000000",
                                952 => "0011001000",
                                953 => "1011000100",
                                954 => "1000110000",
                                955 => "0100011100",
                                956 => "0100111100",
                                957 => "0000100000",
                                958 => "0000000000",
                                959 => "0100010101",
                                960 => "0100010110",
                                961 => "0000000000",
                                962 => "0000000000",
                                963 => "0011000000",
                                964 => "1001110100",
                                965 => "1101111100",
                                966 => "0000000000",
                                967 => "0000000000",
                                968 => "1111001100",
                                969 => "0000011000",
                                970 => "1110010000",
                                971 => "0000001000",
                                972 => "1000111100",
                                973 => "1100110000",
                                974 => "1111010000",
                                975 => "0000101000",
                                976 => "1100000000",
                                977 => "1010100000",
                                978 => "0000000100",
                                979 => "0110011000",
                                980 => "0000000100",
                                981 => "1011101100",
                                982 => "1110010000",
                                983 => "1101010000",
                                984 => "0110100000",
                                985 => "1101111100",
                                986 => "1111001000",
                                987 => "0010110000",
                                988 => "1101110100",
                                989 => "1111010100",
                                990 => "1001011100",
                                991 => "0001100100",
                                992 => "0111000000",
                                993 => "0001001000",
                                994 => "0000010100",
                                995 => "1010000000",
                                996 => "1000000000",
                                997 => "1111001000",
                                998 => "0000000000",
                                999 => "0000000000",
                                1000 => "0000001000",
                                1001 => "0000010000",
                                1002 => "0000010100",
                                1003 => "1010000000",
                                1004 => "0000000100",
                                1005 => "0000000100",
                                1006 => "0000010000",
                                1007 => "0000001000",
                                1008 => "1001110000",
                                1009 => "1011011000",
                                1010 => "1101000000",
                                1011 => "0001011100",
                                1012 => "0100101100",
                                1013 => "0000100100",
                                1014 => "0110000000",
                                1015 => "0011001000",
                                1016 => "1011000100",
                                1017 => "1000110000",
                                1018 => "0100011100",
                                1019 => "0100111100",
                                1020 => "0000100000",
                                1021 => "0000000000",
                                1022 => "0100010101",
                                1023 => "0100010110",
                                1024 => "0000100000",
                                1025 => "0000000000",
                                1026 => "0011000000",
                                1027 => "0101110100",
                                1028 => "1001011000",
                                1029 => "0100000000",
                                1030 => "0000000000",
                                1031 => "0111001100",
                                1032 => "0000011000",
                                1033 => "0110100100",
                                1034 => "1011011100",
                                1035 => "1100011100",
                                1036 => "0100011100",
                                1037 => "1011011100",
                                1038 => "0001110000",
                                1039 => "1100000000",
                                1040 => "1010100000",
                                1041 => "0000000100",
                                1042 => "0110011000",
                                1043 => "0000000100",
                                1044 => "1011101100",
                                1045 => "1110010000",
                                1046 => "1101000000",
                                1047 => "0101010100",
                                1048 => "0101101100",
                                1049 => "1011100100",
                                1050 => "0101111100",
                                1051 => "1111001100",
                                1052 => "0010011100",
                                1053 => "1100010000",
                                1054 => "0100110100",
                                1055 => "0111000000",
                                1056 => "0001001000",
                                1057 => "0010000000",
                                1058 => "0000000000",
                                1059 => "0111010100",
                                1060 => "1110000000",
                                1061 => "0000000000",
                                1062 => "0000000000",
                                1063 => "0000001000",
                                1064 => "0000010000",
                                1065 => "0000010100",
                                1066 => "1011010000",
                                1067 => "0000000100",
                                1068 => "0000000100",
                                1069 => "0000010000",
                                1070 => "0000001000",
                                1071 => "1001110000",
                                1072 => "1011011000",
                                1073 => "1101000000",
                                1074 => "0001011100",
                                1075 => "0100101100",
                                1076 => "0000100100",
                                1077 => "0110000000",
                                1078 => "0011001000",
                                1079 => "1011000100",
                                1080 => "1000110000",
                                1081 => "0100011100",
                                1082 => "0100111100",
                                1083 => "0000100000",
                                1084 => "0000000000",
                                1085 => "0100010101",
                                1086 => "0100010110",
                                1087 => "0000100000",
                                1088 => "0000000000",
                                1089 => "0011000000",
                                1090 => "0101110100",
                                1091 => "1001011100",
                                1092 => "0100000000",
                                1093 => "0000000000",
                                1094 => "0111001100",
                                1095 => "0000011000",
                                1096 => "0110100100",
                                1097 => "1011011000",
                                1098 => "1100011100",
                                1099 => "0100011100",
                                1100 => "1011011100",
                                1101 => "0001110000",
                                1102 => "1100000000",
                                1103 => "1010100000",
                                1104 => "0000000100",
                                1105 => "0110011000",
                                1106 => "0000000100",
                                1107 => "1011101100",
                                1108 => "1110010000",
                                1109 => "1101000100",
                                1110 => "0000101100",
                                1111 => "0010010100",
                                1112 => "1110010000",
                                1113 => "0010100100",
                                1114 => "0110101100",
                                1115 => "0000011100",
                                1116 => "0011000100",
                                1117 => "1011110100",
                                1118 => "0111000000",
                                1119 => "0001001000",
                                1120 => "0010000000",
                                1121 => "0000000000",
                                1122 => "1010111100",
                                1123 => "1111110000",
                                1124 => "0000000000",
                                1125 => "0000000000",
                                1126 => "0000001000",
                                1127 => "0000010000",
                                1128 => "0000010100",
                                1129 => "1011010000",
                                1130 => "0000000100",
                                1131 => "0000000100",
                                1132 => "0000010000",
                                1133 => "0000001000",
                                1134 => "1001110000",
                                1135 => "1011011000",
                                1136 => "1101000000",
                                1137 => "0001011100",
                                1138 => "0100101100",
                                1139 => "0000100100",
                                1140 => "0110000000",
                                1141 => "0011001000",
                                1142 => "1011000100",
                                1143 => "1000110000",
                                1144 => "0100011100",
                                1145 => "0100111100",
                                1146 => "0000100000",
                                1147 => "0000000000",
                                1148 => "0100010101",
                                1149 => "0100010110",
                                1150 => "1000000000",
                                1151 => "0000000000",
                                1152 => "0011000000",
                                1153 => "0000011100",
                                1154 => "0101110000",
                                1155 => "0000000000",
                                1156 => "0000000000",
                                1157 => "0111011100",
                                1158 => "0000011000",
                                1159 => "1011100100",
                                1160 => "1100001000",
                                1161 => "1010110000",
                                1162 => "1101100100",
                                1163 => "0001001100",
                                1164 => "0100001000",
                                1165 => "1100000000",
                                1166 => "1010100000",
                                1167 => "0000000100",
                                1168 => "0110011000",
                                1169 => "0000000100",
                                1170 => "1011101100",
                                1171 => "1110010000",
                                1172 => "1101010100",
                                1173 => "1000110000",
                                1174 => "1100101100",
                                1175 => "0011001000",
                                1176 => "1111010000",
                                1177 => "0101110100",
                                1178 => "1101001000",
                                1179 => "1110000100",
                                1180 => "1011101100",
                                1181 => "0111000000",
                                1182 => "0001001000",
                                1183 => "1111111100",
                                1184 => "1111111100",
                                1185 => "0001101100",
                                1186 => "0010010100",
                                1187 => "0000000000",
                                1188 => "0000000000",
                                1189 => "0000001000",
                                1190 => "0000010000",
                                1191 => "0000010100",
                                1192 => "1001011000",
                                1193 => "0000000100",
                                1194 => "0000000100",
                                1195 => "0000010000",
                                1196 => "0000001000",
                                1197 => "1001110000",
                                1198 => "1011011000",
                                1199 => "1101000000",
                                1200 => "0001011100",
                                1201 => "0100101100",
                                1202 => "0000100100",
                                1203 => "0110000000",
                                1204 => "0011001000",
                                1205 => "1011000100",
                                1206 => "1000110000",
                                1207 => "0100011100",
                                1208 => "0100111100",
                                1209 => "0000100000",
                                1210 => "0000000000",
                                1211 => "0100010101",
                                1212 => "0100010110",
                                1213 => "0000000000",
                                1214 => "0000000000",
                                1215 => "0011000000",
                                1216 => "0000000000",
                                1217 => "0000000000",
                                1218 => "0100000000",
                                1219 => "0000000000",
                                1220 => "1110010100",
                                1221 => "0000011000",
                                1222 => "0110011100",
                                1223 => "1110010100",
                                1224 => "0011011000",
                                1225 => "1010101100",
                                1226 => "0011010100",
                                1227 => "0010100100",
                                1228 => "1100000000",
                                1229 => "1010100000",
                                1230 => "0000000100",
                                1231 => "0110011000",
                                1232 => "0000000100",
                                1233 => "1011101100",
                                1234 => "1110010000",
                                1235 => "1101011000",
                                1236 => "0001110100",
                                1237 => "1000010100",
                                1238 => "1010101100",
                                1239 => "1110001100",
                                1240 => "1000001100",
                                1241 => "0000110000",
                                1242 => "0010010000",
                                1243 => "0111111100",
                                1244 => "0111000000",
                                1245 => "0001001000",
                                1246 => "0110100100",
                                1247 => "0000001100",
                                1248 => "1001010000",
                                1249 => "1010001100",
                                1250 => "0000000000",
                                1251 => "0000000000",
                                1252 => "0000001000",
                                1253 => "0000010000",
                                1254 => "0000010100",
                                1255 => "1011010000",
                                1256 => "0000000100",
                                1257 => "0000000100",
                                1258 => "0000010000",
                                1259 => "0000001000",
                                1260 => "1001110000",
                                1261 => "1011011000",
                                1262 => "1101000000",
                                1263 => "0001011100",
                                1264 => "0100101100",
                                1265 => "0000100100",
                                1266 => "0110000000",
                                1267 => "0011001000",
                                1268 => "1011000100",
                                1269 => "1000110000",
                                1270 => "0100011100",
                                1271 => "0100111100",
                                1272 => "0000100000",
                                1273 => "0000000000",
                                1274 => "0100010101",
                                1275 => "0100010110",
                                1276 => "0000000000",
                                1277 => "0000000000",
                                1278 => "0011000000",
                                1279 => "0000000000",
                                1280 => "0000000000",
                                1281 => "0100000000",
                                1282 => "0000000000",
                                1283 => "1110110000",
                                1284 => "0000011000",
                                1285 => "1111101000",
                                1286 => "0010000100",
                                1287 => "0011011000",
                                1288 => "1010010100",
                                1289 => "1001101100",
                                1290 => "1111001000",
                                1291 => "1100000000",
                                1292 => "1010100000",
                                1293 => "0000000100",
                                1294 => "0110011000",
                                1295 => "0000000100",
                                1296 => "1011101100",
                                1297 => "1110010000",
                                1298 => "1101011100",
                                1299 => "1011010100",
                                1300 => "0110101100",
                                1301 => "0110010000",
                                1302 => "0010110100",
                                1303 => "1101111100",
                                1304 => "1110010100",
                                1305 => "0101110100",
                                1306 => "1110010000",
                                1307 => "0111000000",
                                1308 => "0001001000",
                                1309 => "0110100100",
                                1310 => "0000001100",
                                1311 => "0100011100",
                                1312 => "0111000000",
                                1313 => "0000000000",
                                1314 => "0000000000",
                                1315 => "0000001000",
                                1316 => "0000010000",
                                1317 => "0000010100",
                                1318 => "1011010000",
                                1319 => "0000000100",
                                1320 => "0000000100",
                                1321 => "0000010000",
                                1322 => "0000001000",
                                1323 => "1001110000",
                                1324 => "1011011000",
                                1325 => "1101000000",
                                1326 => "0001011100",
                                1327 => "0100101100",
                                1328 => "0000100100",
                                1329 => "0110000000",
                                1330 => "0011001000",
                                1331 => "1011000100",
                                1332 => "1000110000",
                                1333 => "0100011100",
                                1334 => "0100111100",
                                1335 => "0000100000",
                                1336 => "0000000000",
                                1337 => "0100010101",
                                1338 => "0100010110",
                                1339 => "0000000000",
                                1340 => "0000000000",
                                1341 => "0011000000",
                                1342 => "0000000000",
                                1343 => "0000000000",
                                1344 => "0100000000",
                                1345 => "0000000000",
                                1346 => "1110110000",
                                1347 => "0000011000",
                                1348 => "0010111000",
                                1349 => "1001100100",
                                1350 => "0010001100",
                                1351 => "1010110000",
                                1352 => "0111101000",
                                1353 => "0111010000",
                                1354 => "1100000000",
                                1355 => "1010100000",
                                1356 => "0000000100",
                                1357 => "0110011000",
                                1358 => "0000000100",
                                1359 => "1011101100",
                                1360 => "1110010000",
                                1361 => "1101100000",
                                1362 => "1110000000",
                                1363 => "0111110000",
                                1364 => "1011101100",
                                1365 => "1100010100",
                                1366 => "1100010100",
                                1367 => "0000110100",
                                1368 => "0001001100",
                                1369 => "0010110100",
                                1370 => "0111000000",
                                1371 => "0001001000",
                                1372 => "0110100100",
                                1373 => "0000001100",
                                1374 => "0101111000",
                                1375 => "1100110000",
                                1376 => "0000000000",
                                1377 => "0000000000",
                                1378 => "0000001000",
                                1379 => "0000010000",
                                1380 => "0000010100",
                                1381 => "1011010000",
                                1382 => "0000000100",
                                1383 => "0000000100",
                                1384 => "0000010000",
                                1385 => "0000001000",
                                1386 => "1001110000",
                                1387 => "1011011000",
                                1388 => "1101000000",
                                1389 => "0001011100",
                                1390 => "0100101100",
                                1391 => "0000100100",
                                1392 => "0110000000",
                                1393 => "0011001000",
                                1394 => "1011000100",
                                1395 => "1000110000",
                                1396 => "0100011100",
                                1397 => "0100111100",
                                1398 => "0000100000",
                                1399 => "0000000000",
                                1400 => "0100010101",
                                1401 => "0100010110",
                                1402 => "0000000000",
                                1403 => "0000000000",
                                1404 => "0011000000",
                                1405 => "0000000000",
                                1406 => "0000000000",
                                1407 => "0100000000",
                                1408 => "0000000000",
                                1409 => "0011000100",
                                1410 => "0000011000",
                                1411 => "0111110100",
                                1412 => "1001101000",
                                1413 => "1011100100",
                                1414 => "1001111100",
                                1415 => "0101000000",
                                1416 => "1000000000",
                                1417 => "1100000000",
                                1418 => "1010100000",
                                1419 => "0000000100",
                                1420 => "0110011000",
                                1421 => "0001111100",
                                1422 => "1001110000",
                                1423 => "1110010000",
                                1424 => "1101100100",
                                1425 => "1100000100",
                                1426 => "0010110100",
                                1427 => "1110010000",
                                1428 => "1101001000",
                                1429 => "0111111100",
                                1430 => "0110010000",
                                1431 => "0001101100",
                                1432 => "1111111000",
                                1433 => "0111000000",
                                1434 => "0001001000",
                                1435 => "1010010100",
                                1436 => "0110010000",
                                1437 => "1100101100",
                                1438 => "1010001100",
                                1439 => "0000000000",
                                1440 => "0000000000",
                                1441 => "0000001000",
                                1442 => "0000010000",
                                1443 => "0000010100",
                                1444 => "1011010000",
                                1445 => "0000000100",
                                1446 => "0000000100",
                                1447 => "0000010000",
                                1448 => "0000001000",
                                1449 => "1001110000",
                                1450 => "1011011000",
                                1451 => "1101000000",
                                1452 => "0001011100",
                                1453 => "0100101100",
                                1454 => "0000100100",
                                1455 => "0110000000",
                                1456 => "0011001000",
                                1457 => "1011000100",
                                1458 => "1000110000",
                                1459 => "0100011100",
                                1460 => "0100111100",
                                1461 => "0000100000",
                                1462 => "0000000000",
                                1463 => "0100010101",
                                1464 => "0100010110",
                                1465 => "0000000000",
                                1466 => "0000000000",
                                1467 => "0011000000",
                                1468 => "1100000000",
                                1469 => "1000000100",
                                1470 => "0100000000",
                                1471 => "0000000000",
                                1472 => "0111011100",
                                1473 => "0000011000",
                                1474 => "0101111000",
                                1475 => "0000010100",
                                1476 => "0000110100",
                                1477 => "0110101100",
                                1478 => "0001010100",
                                1479 => "1100100000",
                                1480 => "1100000000",
                                1481 => "1010100000",
                                1482 => "0000000100",
                                1483 => "0110011000",
                                1484 => "0000000100",
                                1485 => "1011101100",
                                1486 => "1110010000",
                                1487 => "1101101000",
                                1488 => "1001011000",
                                1489 => "1010010100",
                                1490 => "0111001100",
                                1491 => "1000101000",
                                1492 => "0000000000",
                                1493 => "1110110000",
                                1494 => "1110110000",
                                1495 => "0010101000",
                                1496 => "0111000000",
                                1497 => "0001001000",
                                1498 => "1111101000",
                                1499 => "1111000000",
                                1500 => "1100010100",
                                1501 => "0001010000",
                                1502 => "0000000000",
                                1503 => "0000000000",
                                1504 => "0000001000",
                                1505 => "0000010000",
                                1506 => "0000010100",
                                1507 => "1010000000",
                                1508 => "0000000100",
                                1509 => "0000000100",
                                1510 => "0000010000",
                                1511 => "0000001000",
                                1512 => "1001110000",
                                1513 => "1011011000",
                                1514 => "1101000000",
                                1515 => "0001011100",
                                1516 => "0100101100",
                                1517 => "0000100100",
                                1518 => "0110000000",
                                1519 => "0011001000",
                                1520 => "1011000100",
                                1521 => "1000110000",
                                1522 => "0100011100",
                                1523 => "0100111100",
                                1524 => "0000100000",
                                1525 => "0000000000",
                                1526 => "0100010101",
                                1527 => "0100010110",
                                1528 => "0000000000",
                                1529 => "0000000000",
                                1530 => "0011000000",
                                1531 => "0000000000",
                                1532 => "0000000000",
                                1533 => "0100000000",
                                1534 => "0000000000",
                                1535 => "0011100000",
                                1536 => "0000011000",
                                1537 => "0010101100",
                                1538 => "0001011100",
                                1539 => "0110100000",
                                1540 => "0111100100",
                                1541 => "1110110100",
                                1542 => "0010100100",
                                1543 => "1100000000",
                                1544 => "1010100000",
                                1545 => "0000000100",
                                1546 => "0110011000",
                                1547 => "0000000100",
                                1548 => "1011101100",
                                1549 => "1110010000",
                                1550 => "1101101100",
                                1551 => "0010010100",
                                1552 => "1000101000",
                                1553 => "1010110100",
                                1554 => "0000000000",
                                1555 => "0000101000",
                                1556 => "0011010100",
                                1557 => "1111000000",
                                1558 => "1101011100",
                                1559 => "0111000000",
                                1560 => "0001001000",
                                1561 => "1111101000",
                                1562 => "1111000000",
                                1563 => "1011110000",
                                1564 => "0011111000",
                                1565 => "0000000000",
                                1566 => "0000000000",
                                1567 => "0000001000",
                                1568 => "0000010000",
                                1569 => "0000010100",
                                1570 => "1011010000",
                                1571 => "0000000100",
                                1572 => "0000000100",
                                1573 => "0000010000",
                                1574 => "0000001000",
                                1575 => "1001110000",
                                1576 => "1011011000",
                                1577 => "1101000000",
                                1578 => "0001011100",
                                1579 => "0100101100",
                                1580 => "0000100100",
                                1581 => "0110000000",
                                1582 => "0011001000",
                                1583 => "1011000100",
                                1584 => "1000110000",
                                1585 => "0100011100",
                                1586 => "0100111100",
                                1587 => "0000100000",
                                1588 => "0000000000",
                                1589 => "0100010101",
                                1590 => "0100010110",
                                1591 => "0000000000",
                                1592 => "0000000000",
                                1593 => "0011000000",
                                1594 => "0000000000",
                                1595 => "0000000000",
                                1596 => "0100000000",
                                1597 => "0000000000",
                                1598 => "0011011000",
                                1599 => "0000011000",
                                1600 => "1001001000",
                                1601 => "1001101000",
                                1602 => "0000001000",
                                1603 => "0001011000",
                                1604 => "1110111000",
                                1605 => "0000100100",
                                1606 => "1100000000",
                                1607 => "1010100000",
                                1608 => "0000000100",
                                1609 => "0110011000",
                                1610 => "0000000100",
                                1611 => "1011101100",
                                1612 => "1110010000",
                                1613 => "1101110000",
                                1614 => "0100100100",
                                1615 => "0110010100",
                                1616 => "0101011100",
                                1617 => "1110111100",
                                1618 => "0101001000",
                                1619 => "0111100000",
                                1620 => "0001000100",
                                1621 => "1101010100",
                                1622 => "0111000000",
                                1623 => "0001001000",
                                1624 => "1111101000",
                                1625 => "1111000000",
                                1626 => "1110100100",
                                1627 => "1011011000",
                                1628 => "0000000000",
                                1629 => "0000000000",
                                1630 => "0000001000",
                                1631 => "0000010000",
                                1632 => "0000010100",
                                1633 => "1011010000",
                                1634 => "0000000100",
                                1635 => "0000000100",
                                1636 => "0000010000",
                                1637 => "0000001000",
                                1638 => "1001110000",
                                1639 => "1011011000",
                                1640 => "1101000000",
                                1641 => "0001011100",
                                1642 => "0100101100",
                                1643 => "0000100100",
                                1644 => "0110000000",
                                1645 => "0011001000",
                                1646 => "1011000100",
                                1647 => "1000110000",
                                1648 => "0100011100",
                                1649 => "0100111100",
                                1650 => "0000100000",
                                1651 => "0000000000",
                                1652 => "0100010101",
                                1653 => "0100010110",
                                1654 => "0000000000",
                                1655 => "0000000000",
                                1656 => "0011000000",
                                1657 => "0000000000",
                                1658 => "0000000000",
                                1659 => "0100000000",
                                1660 => "0000000000",
                                1661 => "0011011000",
                                1662 => "0000011000",
                                1663 => "1001001000",
                                1664 => "1001101000",
                                1665 => "0000001000",
                                1666 => "0001011000",
                                1667 => "1110111000",
                                1668 => "0000100100",
                                1669 => "1100000000",
                                1670 => "1010100000",
                                1671 => "0000000100",
                                1672 => "0110011000",
                                1673 => "0000000100",
                                1674 => "1011101100",
                                1675 => "1110010000",
                                1676 => "1101111000",
                                1677 => "1101000100",
                                1678 => "1001110000",
                                1679 => "1011001000",
                                1680 => "1100010100",
                                1681 => "1101110100",
                                1682 => "0010100000",
                                1683 => "1011011100",
                                1684 => "0000101000",
                                1685 => "0111000000",
                                1686 => "0001001000",
                                1687 => "1111101000",
                                1688 => "1111000000",
                                1689 => "1101011000",
                                1690 => "1100000000",
                                1691 => "0000000000",
                                1692 => "0000000000",
                                1693 => "0000001000",
                                1694 => "0000010000",
                                1695 => "0000010100",
                                1696 => "1011010000",
                                1697 => "0000000100",
                                1698 => "0000000100",
                                1699 => "0000010000",
                                1700 => "0000001000",
                                1701 => "1001110000",
                                1702 => "1011011000",
                                1703 => "1101000000",
                                1704 => "0001011100",
                                1705 => "0100101100",
                                1706 => "0000100100",
                                1707 => "0110000000",
                                1708 => "0011001000",
                                1709 => "1011000100",
                                1710 => "1000110000",
                                1711 => "0100011100",
                                1712 => "0100111100",
                                1713 => "0000100000",
                                1714 => "0000000000",
                                1715 => "0100010101",
                                1716 => "0100010110",
                                1717 => "0000000000",
                                1718 => "0000000000",
                                1719 => "0011000000",
                                1720 => "0000000000",
                                1721 => "0000000000",
                                1722 => "0100000000",
                                1723 => "0000000000",
                                1724 => "1110110000",
                                1725 => "0000011000",
                                1726 => "0010111000",
                                1727 => "1001100100",
                                1728 => "0010001100",
                                1729 => "1010110000",
                                1730 => "0111101000",
                                1731 => "0111010000",
                                1732 => "1100000000",
                                1733 => "1010100000",
                                1734 => "0000000100",
                                1735 => "0110011000",
                                1736 => "0000000100",
                                1737 => "1011101100",
                                1738 => "1110010000",
                                1739 => "1101110100",
                                1740 => "0111111000",
                                1741 => "1100110100",
                                1742 => "0100100100",
                                1743 => "1100101000",
                                1744 => "1010100100",
                                1745 => "1000111000",
                                1746 => "1100000000",
                                1747 => "1000011100",
                                1748 => "0111000000",
                                1749 => "0001001000",
                                1750 => "0110100100",
                                1751 => "0000001100",
                                1752 => "1010000000",
                                1753 => "1001011000",
                                1754 => "0000000000",
                                1755 => "0000000000",
                                1756 => "0000001000",
                                1757 => "0000010000",
                                1758 => "0000010100",
                                1759 => "1011010000",
                                1760 => "0000000100",
                                1761 => "0000000100",
                                1762 => "0000010000",
                                1763 => "0000001000",
                                1764 => "1001110000",
                                1765 => "1011011000",
                                1766 => "1101000000",
                                1767 => "0001011100",
                                1768 => "0100101100",
                                1769 => "0000100100",
                                1770 => "0110000000",
                                1771 => "0011001000",
                                1772 => "1011000100",
                                1773 => "1000110000",
                                1774 => "0100011100",
                                1775 => "0100111100",
                                1776 => "0000100000",
                                1777 => "0000000000",
                                1778 => "0100010101",
                                1779 => "0100010110",
                                1780 => "0000000000",
                                1781 => "0000000000",
                                1782 => "0011000000",
                                1783 => "0000000000",
                                1784 => "0000000000",
                                1785 => "0100000000",
                                1786 => "0000000000",
                                1787 => "1110010000",
                                1788 => "0000011000",
                                1789 => "0111000100",
                                1790 => "1101110000",
                                1791 => "0011111100",
                                1792 => "0010000100",
                                1793 => "0010001100",
                                1794 => "1011110000",
                                1795 => "1100000000",
                                1796 => "1010100000",
                                1797 => "0000000100",
                                1798 => "0110011000",
                                1799 => "0000000100",
                                1800 => "1011101100",
                                1801 => "1110010000",
                                1802 => "1101111100",
                                1803 => "1111110100",
                                1804 => "0111110100",
                                1805 => "1101101000",
                                1806 => "0100010100",
                                1807 => "0110110100",
                                1808 => "0000000100",
                                1809 => "1000001000",
                                1810 => "0101000100",
                                1811 => "0111000000",
                                1812 => "0001001000",
                                1813 => "0110100100",
                                1814 => "0000001100",
                                1815 => "0100011100",
                                1816 => "0110111100",
                                1817 => "0000000000",
                                1818 => "0000000000",
                                1819 => "0000001000",
                                1820 => "0000010000",
                                1821 => "0000010100",
                                1822 => "1011010000",
                                1823 => "0000000100",
                                1824 => "0000000100",
                                1825 => "0000010000",
                                1826 => "0000001000",
                                1827 => "1001110000",
                                1828 => "1011011000",
                                1829 => "1101000000",
                                1830 => "0001011100",
                                1831 => "0100101100",
                                1832 => "0000100100",
                                1833 => "0110000000",
                                1834 => "0011001000",
                                1835 => "1011000100",
                                1836 => "1000110000",
                                1837 => "0100011100",
                                1838 => "0100111100",
                                1839 => "0000100000",
                                1840 => "0000000000",
                                1841 => "0100010101",
                                1842 => "0100010110",
                                1843 => "0000000000",
                                1844 => "0000000000",
                                1845 => "0011000000",
                                1846 => "0000000000",
                                1847 => "0000000000",
                                1848 => "0100000000",
                                1849 => "0000000000",
                                1850 => "0011100100",
                                1851 => "0000011000",
                                1852 => "0111001000",
                                1853 => "1001000100",
                                1854 => "1100000000",
                                1855 => "0000000000",
                                1856 => "0100110100",
                                1857 => "0010100000",
                                1858 => "1100000000",
                                1859 => "1010100000",
                                1860 => "0000000100",
                                1861 => "0110011000",
                                1862 => "0000000100",
                                1863 => "1011101100",
                                1864 => "1110010000",
                                1865 => "1110000000",
                                1866 => "1001101100",
                                1867 => "1100001000",
                                1868 => "0110001000",
                                1869 => "1000011100",
                                1870 => "1000001000",
                                1871 => "1101000100",
                                1872 => "0100100100",
                                1873 => "1101111000",
                                1874 => "0111000000",
                                1875 => "0001001000",
                                1876 => "0111001000",
                                1877 => "0001000000",
                                1878 => "1001000000",
                                1879 => "0011001000",
                                1880 => "0000000000",
                                1881 => "0000000000",
                                1882 => "0000001000",
                                1883 => "0000010000",
                                1884 => "0000010100",
                                1885 => "1011010000",
                                1886 => "0000000100",
                                1887 => "0000000100",
                                1888 => "0000010000",
                                1889 => "0000001000",
                                1890 => "1001110000",
                                1891 => "1011011000",
                                1892 => "1101000000",
                                1893 => "0001011100",
                                1894 => "0100101100",
                                1895 => "0000100100",
                                1896 => "0110000000",
                                1897 => "0011001000",
                                1898 => "1011000100",
                                1899 => "1000110000",
                                1900 => "0100011100",
                                1901 => "0100111100",
                                1902 => "0000100000",
                                1903 => "0000000000",
                                1904 => "0100010101",
                                1905 => "0100010110",
                                1906 => "0000000000",
                                1907 => "0000000000",
                                1908 => "0011000000",
                                1909 => "1001010100",
                                1910 => "0001001000",
                                1911 => "0000000000",
                                1912 => "0000000000",
                                1913 => "1111001100",
                                1914 => "0000011000",
                                1915 => "1100101100",
                                1916 => "0011110100",
                                1917 => "0000110100",
                                1918 => "0010000100",
                                1919 => "1001100000",
                                1920 => "0100100000",
                                1921 => "1100000000",
                                1922 => "1010100000",
                                1923 => "0000000100",
                                1924 => "0110011000",
                                1925 => "0000000100",
                                1926 => "1011101100",
                                1927 => "1110010000",
                                1928 => "1110000100",
                                1929 => "0100101000",
                                1930 => "0001001100",
                                1931 => "1110010100",
                                1932 => "0100001000",
                                1933 => "1001001100",
                                1934 => "1100011000",
                                1935 => "1111101100",
                                1936 => "0000100000",
                                1937 => "0111000000",
                                1938 => "0001001000",
                                1939 => "0000010100",
                                1940 => "1010000000",
                                1941 => "0111000100",
                                1942 => "0100100100",
                                1943 => "0000000000",
                                1944 => "0000000000",
                                1945 => "0000001000",
                                1946 => "0000010000",
                                1947 => "0000010100",
                                1948 => "1010000000",
                                1949 => "0000000100",
                                1950 => "0000000100",
                                1951 => "0000010000",
                                1952 => "0000001000",
                                1953 => "1001110000",
                                1954 => "1011011000",
                                1955 => "1101000000",
                                1956 => "0001011100",
                                1957 => "0100101100",
                                1958 => "0000100100",
                                1959 => "0110000000",
                                1960 => "0011001000",
                                1961 => "1011000100",
                                1962 => "1000110000",
                                1963 => "0100011100",
                                1964 => "0100111100",
                                1965 => "0000100000",
                                1966 => "0000000000",
                                1967 => "0100010101",
                                1968 => "0100010110",
                                1969 => "0000000000",
                                1970 => "0000000000",
                                1971 => "0011000000",
                                1972 => "1110001000",
                                1973 => "1100001100",
                                1974 => "0100000000",
                                1975 => "0000000000",
                                1976 => "0011010100",
                                1977 => "0000011000",
                                1978 => "0001011000",
                                1979 => "1001010000",
                                1980 => "0100010100",
                                1981 => "0101101000",
                                1982 => "0100010100",
                                1983 => "0000100000",
                                1984 => "1100000000",
                                1985 => "1010100000",
                                1986 => "0000000100",
                                1987 => "0110011000",
                                1988 => "0000000100",
                                1989 => "1011101100",
                                1990 => "1110010000",
                                1991 => "1110001000",
                                1992 => "0101110000",
                                1993 => "0101101100",
                                1994 => "0110111100",
                                1995 => "1000001100",
                                1996 => "1011110100",
                                1997 => "1001001100",
                                1998 => "1101011000",
                                1999 => "1100100000",
                                2000 => "0111000000",
                                2001 => "0001001000",
                                2002 => "0001011000",
                                2003 => "1101000000",
                                2004 => "1101100000",
                                2005 => "1111010100",
                                2006 => "0000000000",
                                2007 => "0000000000",
                                2008 => "0000001000",
                                2009 => "0000010000",
                                2010 => "0000010100",
                                2011 => "1011010000",
                                2012 => "0000000100",
                                2013 => "0000000100",
                                2014 => "0000010000",
                                2015 => "0000001000",
                                2016 => "1001110000",
                                2017 => "1011011000",
                                2018 => "1101000000",
                                2019 => "0001011100",
                                2020 => "0100101100",
                                2021 => "0000100100",
                                2022 => "0110000000",
                                2023 => "0011001000",
                                2024 => "1011000100",
                                2025 => "1000110000",
                                2026 => "0100011100",
                                2027 => "0100111100",
                                2028 => "0000100000",
                                2029 => "0000000000",
                                2030 => "0100010101",
                                2031 => "0100010110",
                                2032 => "0000000000",
                                2033 => "0000000000",
                                2034 => "0011000000",
                                2035 => "1110010000",
                                2036 => "1100001100",
                                2037 => "0100000000",
                                2038 => "0000000000",
                                2039 => "0011010100",
                                2040 => "0000011000",
                                2041 => "0001010000",
                                2042 => "1001010000",
                                2043 => "0100010100",
                                2044 => "0101101000",
                                2045 => "0100010100",
                                2046 => "0000100000",
                                2047 => "1100000000",
                                2048 => "1010100000",
                                2049 => "0000000100",
                                2050 => "0110011000",
                                2051 => "0000000100",
                                2052 => "1011101100",
                                2053 => "1110010000",
                                2054 => "1110001100",
                                2055 => "0111001100",
                                2056 => "0111001000",
                                2057 => "0111001100",
                                2058 => "1101100100",
                                2059 => "1111001000",
                                2060 => "0100001000",
                                2061 => "0110111100",
                                2062 => "0101101000",
                                2063 => "0111000000",
                                2064 => "0001001000",
                                2065 => "0001011000",
                                2066 => "1101000000",
                                2067 => "1111000000",
                                2068 => "0100011000",
                                2069 => "0000000000",
                                2070 => "0000000000",
                                2071 => "0000001000",
                                2072 => "0000010000",
                                2073 => "0000010100",
                                2074 => "1011010000",
                                2075 => "0000000100",
                                2076 => "0000000100",
                                2077 => "0000010000",
                                2078 => "0000001000",
                                2079 => "1001110000",
                                2080 => "1011011000",
                                2081 => "1101000000",
                                2082 => "0001011100",
                                2083 => "0100101100",
                                2084 => "0000100100",
                                2085 => "0110000000",
                                2086 => "0011001000",
                                2087 => "1011000100",
                                2088 => "1000110000",
                                2089 => "0100011100",
                                2090 => "0100111100",
                                2091 => "0000100000",
                                2092 => "0000000000",
                                2093 => "0100010101",
                                2094 => "0100010110",
                                2095 => "0000000000",
                                2096 => "0000000000",
                                2097 => "0011000000",
                                2098 => "0000000000",
                                2099 => "0000000000",
                                2100 => "0100000000",
                                2101 => "0000000000",
                                2102 => "0011100100",
                                2103 => "0000011000",
                                2104 => "0111001100",
                                2105 => "1011011000",
                                2106 => "1100000000",
                                2107 => "0000000000",
                                2108 => "0100110000",
                                2109 => "0000001100",
                                2110 => "1100000000",
                                2111 => "1010100000",
                                2112 => "0000000100",
                                2113 => "0110011000",
                                2114 => "0000000100",
                                2115 => "1011101100",
                                2116 => "1110010000",
                                2117 => "1110010000",
                                2118 => "1010101100",
                                2119 => "1011001100",
                                2120 => "1010000000",
                                2121 => "0001101100",
                                2122 => "1001111000",
                                2123 => "1011001100",
                                2124 => "1101011100",
                                2125 => "1000010100",
                                2126 => "0111000000",
                                2127 => "0001001000",
                                2128 => "0111001000",
                                2129 => "0001000000",
                                2130 => "1001101000",
                                2131 => "0100010000",
                                2132 => "0000000000",
                                2133 => "0000000000",
                                2134 => "0000001000",
                                2135 => "0000010000",
                                2136 => "0000010100",
                                2137 => "1011010000",
                                2138 => "0000000100",
                                2139 => "0000000100",
                                2140 => "0000010000",
                                2141 => "0000001000",
                                2142 => "1001110000",
                                2143 => "1011011000",
                                2144 => "1101000000",
                                2145 => "0001011100",
                                2146 => "0100101100",
                                2147 => "0000100100",
                                2148 => "0110000000",
                                2149 => "0011001000",
                                2150 => "1011000100",
                                2151 => "1000110000",
                                2152 => "0100011100",
                                2153 => "0100111100",
                                2154 => "0000100000",
                                2155 => "0000000000",
                                2156 => "0100010101",
                                2157 => "0100010110",
                                2158 => "0000000000",
                                2159 => "0000000000",
                                2160 => "0011000000",
                                2161 => "0000000000",
                                2162 => "0000000000",
                                2163 => "0100000000",
                                2164 => "0000000000",
                                2165 => "0011100100",
                                2166 => "0000011000",
                                2167 => "0011010100",
                                2168 => "1000110000",
                                2169 => "0001011100",
                                2170 => "1100100100",
                                2171 => "0011001000",
                                2172 => "0110010100",
                                2173 => "1100000000",
                                2174 => "1010100000",
                                2175 => "0000000100",
                                2176 => "0110011000",
                                2177 => "0000000100",
                                2178 => "1011101100",
                                2179 => "1110010000",
                                2180 => "1110010100",
                                2181 => "0111100100",
                                2182 => "0000101100",
                                2183 => "0001101000",
                                2184 => "1011110100",
                                2185 => "1011101000",
                                2186 => "1000010100",
                                2187 => "0100010100",
                                2188 => "1011011100",
                                2189 => "0111000000",
                                2190 => "0001001000",
                                2191 => "1111101000",
                                2192 => "1111000000",
                                2193 => "0000000100",
                                2194 => "0011110000",
                                2195 => "0000000000",
                                2196 => "0000000000",
                                2197 => "0000001000",
                                2198 => "0000010000",
                                2199 => "0000010100",
                                2200 => "1011010000",
                                2201 => "0000000100",
                                2202 => "0000000100",
                                2203 => "0000010000",
                                2204 => "0000001000",
                                2205 => "1001110000",
                                2206 => "1011011000",
                                2207 => "1101000000",
                                2208 => "0001011100",
                                2209 => "0100101100",
                                2210 => "0000100100",
                                2211 => "0110000000",
                                2212 => "0011001000",
                                2213 => "1011000100",
                                2214 => "1000110000",
                                2215 => "0100011100",
                                2216 => "0100111100",
                                2217 => "0000100000",
                                2218 => "0000000000",
                                2219 => "0100010101",
                                2220 => "0100010110",
                                2221 => "0000000000",
                                2222 => "0000000000",
                                2223 => "0011000000",
                                2224 => "0000000000",
                                2225 => "0000000000",
                                2226 => "0100000000",
                                2227 => "0000000000",
                                2228 => "0010100100",
                                2229 => "0000011000",
                                2230 => "0010000000",
                                2231 => "0001100100",
                                2232 => "0000111100",
                                2233 => "1011110000",
                                2234 => "0101111100",
                                2235 => "1110010100",
                                2236 => "1100000000",
                                2237 => "1010100000",
                                2238 => "0000000100",
                                2239 => "0110011000",
                                2240 => "0000000100",
                                2241 => "1011101100",
                                2242 => "1110010000",
                                2243 => "1110011000",
                                2244 => "1100001100",
                                2245 => "0111010000",
                                2246 => "0111110000",
                                2247 => "1110101100",
                                2248 => "0100001100",
                                2249 => "1001000100",
                                2250 => "1110011000",
                                2251 => "1111011000",
                                2252 => "0111000000",
                                2253 => "0001001000",
                                2254 => "1111111100",
                                2255 => "1111111100",
                                2256 => "1111111100",
                                2257 => "1101010100",
                                2258 => "0000000000",
                                2259 => "0000000000",
                                2260 => "0000001000",
                                2261 => "0000010000",
                                2262 => "0000010100",
                                2263 => "1011010000",
                                2264 => "0000000100",
                                2265 => "0000000100",
                                2266 => "0000010000",
                                2267 => "0000001000",
                                2268 => "1001110000",
                                2269 => "1011011000",
                                2270 => "1101000000",
                                2271 => "0001011100",
                                2272 => "0100101100",
                                2273 => "0000100100",
                                2274 => "0110000000",
                                2275 => "0011001000",
                                2276 => "1011000100",
                                2277 => "1000110000",
                                2278 => "0100011100",
                                2279 => "0100111100",
                                2280 => "0000100000",
                                2281 => "0000000000",
                                2282 => "0100010101",
                                2283 => "0100010110",
                                2284 => "0000000000",
                                2285 => "0000000000",
                                2286 => "0011000000",
                                2287 => "1011000000",
                                2288 => "0011001000",
                                2289 => "0000000000",
                                2290 => "0000000000",
                                2291 => "1111010000",
                                2292 => "0000011000",
                                2293 => "1101000000",
                                2294 => "1010111100",
                                2295 => "1000111100",
                                2296 => "1100110000",
                                2297 => "1111010000",
                                2298 => "0000101000",
                                2299 => "1100000000",
                                2300 => "1010100000",
                                2301 => "0000000100",
                                2302 => "0110011000",
                                2303 => "0000000100",
                                2304 => "1011101100",
                                2305 => "1110010000",
                                2306 => "1110011100",
                                2307 => "0011010000",
                                2308 => "0000111000",
                                2309 => "1100001000",
                                2310 => "0010001100",
                                2311 => "0011101100",
                                2312 => "0100100000",
                                2313 => "0101011100",
                                2314 => "0110001000",
                                2315 => "0111000000",
                                2316 => "0001001000",
                                2317 => "0000010100",
                                2318 => "1010000000",
                                2319 => "1100100000",
                                2320 => "0001111000",
                                2321 => "0000000000",
                                2322 => "0000000000",
                                2323 => "0000001000",
                                2324 => "0000010000",
                                2325 => "0000010100",
                                2326 => "1010000000",
                                2327 => "0000000100",
                                2328 => "0000000100",
                                2329 => "0000010000",
                                2330 => "0000001000",
                                2331 => "1001110000",
                                2332 => "1011011000",
                                2333 => "1101000000",
                                2334 => "0001011100",
                                2335 => "0100101100",
                                2336 => "0000100100",
                                2337 => "0110000000",
                                2338 => "0011001000",
                                2339 => "1011000100",
                                2340 => "1000110000",
                                2341 => "0100011100",
                                2342 => "0100111100",
                                2343 => "0000100000",
                                2344 => "0000000000",
                                2345 => "0100010101",
                                2346 => "0100010110",
                                2347 => "0000000000",
                                2348 => "0000000000",
                                2349 => "0011000000",
                                2350 => "1010001000",
                                2351 => "0010000100",
                                2352 => "0100000000",
                                2353 => "0000000000",
                                2354 => "0111011000",
                                2355 => "0000011000",
                                2356 => "0110100100",
                                2357 => "0001111100",
                                2358 => "0000110100",
                                2359 => "0110101100",
                                2360 => "0010101000",
                                2361 => "0000111000",
                                2362 => "1100000000",
                                2363 => "1010100000",
                                2364 => "0000000100",
                                2365 => "0110011000",
                                2366 => "0000000100",
                                2367 => "1011101100",
                                2368 => "1110010000",
                                2369 => "1110100000",
                                2370 => "1000111100",
                                2371 => "0010010000",
                                2372 => "0001011000",
                                2373 => "0100100100",
                                2374 => "1110001000",
                                2375 => "1011001000",
                                2376 => "0100000000",
                                2377 => "1110100100",
                                2378 => "0111000000",
                                2379 => "0001001000",
                                2380 => "1111101000",
                                2381 => "1111000000",
                                2382 => "1101111000",
                                2383 => "1111110100",
                                2384 => "0000000000",
                                2385 => "0000000000",
                                2386 => "0000001000",
                                2387 => "0000010000",
                                2388 => "0000010100",
                                2389 => "1010000000",
                                2390 => "0000000100",
                                2391 => "0000000100",
                                2392 => "0000010000",
                                2393 => "0000001000",
                                2394 => "1001110000",
                                2395 => "1011011000",
                                2396 => "1101000000",
                                2397 => "0001011100",
                                2398 => "0100101100",
                                2399 => "0000100100",
                                2400 => "0110000000",
                                2401 => "0011001000",
                                2402 => "1011000100",
                                2403 => "1000110000",
                                2404 => "0100011100",
                                2405 => "0100111100",
                                2406 => "0000100000",
                                2407 => "0000000000",
                                2408 => "0100010101",
                                2409 => "0100010110",
                                2410 => "1000000000",
                                2411 => "0000000000",
                                2412 => "0011000000",
                                2413 => "1111111100",
                                2414 => "1110001000",
                                2415 => "0000000000",
                                2416 => "0000000000",
                                2417 => "0111011100",
                                2418 => "0000011000",
                                2419 => "1010111100",
                                2420 => "0001111000",
                                2421 => "0010001100",
                                2422 => "1111010000",
                                2423 => "1010111000",
                                2424 => "0100010000",
                                2425 => "1100000000",
                                2426 => "1010100000",
                                2427 => "0000000100",
                                2428 => "0110011000",
                                2429 => "0000000100",
                                2430 => "1011101100",
                                2431 => "1110010000",
                                2432 => "1110101000",
                                2433 => "1000100100",
                                2434 => "0110000000",
                                2435 => "1001001100",
                                2436 => "1101000100",
                                2437 => "0010100000",
                                2438 => "0001111100",
                                2439 => "1100110100",
                                2440 => "0000001100",
                                2441 => "0111000000",
                                2442 => "0001001000",
                                2443 => "1111111100",
                                2444 => "1111111100",
                                2445 => "1111010100",
                                2446 => "1110101100",
                                2447 => "0000000000",
                                2448 => "0000000000",
                                2449 => "0000001000",
                                2450 => "0000010000",
                                2451 => "0000010100",
                                2452 => "1001011000",
                                2453 => "0000000100",
                                2454 => "0000000100",
                                2455 => "0000010000",
                                2456 => "0000001000",
                                2457 => "1001110000",
                                2458 => "1011011000",
                                2459 => "1101000000",
                                2460 => "0001011100",
                                2461 => "0100101100",
                                2462 => "0000100100",
                                2463 => "0110000000",
                                2464 => "0011001000",
                                2465 => "1011000100",
                                2466 => "1000110000",
                                2467 => "0100011100",
                                2468 => "0100111100",
                                2469 => "0000100000",
                                2470 => "0000000000",
                                2471 => "0100010101",
                                2472 => "0100010110",
                                2473 => "0000000000",
                                2474 => "0000000000",
                                2475 => "0010110000",
                                2476 => "0000000000",
                                2477 => "0000000000",
                                2478 => "0100000000",
                                2479 => "0000000000",
                                2480 => "1110000100",
                                2481 => "0000011000",
                                2482 => "1001111000",
                                2483 => "0111001100",
                                2484 => "0011011000",
                                2485 => "1110010100",
                                2486 => "0000001000",
                                2487 => "0110010100",
                                2488 => "1100000000",
                                2489 => "1010100000",
                                2490 => "0000000100",
                                2491 => "0110011000",
                                2492 => "0000000100",
                                2493 => "1011101100",
                                2494 => "1110010000",
                                2495 => "1110100100",
                                2496 => "0001011000",
                                2497 => "0101101000",
                                2498 => "0111011000",
                                2499 => "0101111000",
                                2500 => "1001111100",
                                2501 => "0010001100",
                                2502 => "0111000100",
                                2503 => "1001011000",
                                2504 => "0110000000",
                                2505 => "0001001000",
                                2506 => "0110100100",
                                2507 => "0000001100",
                                2508 => "1010111100",
                                2509 => "1010001100",
                                2510 => "0000000000",
                                2511 => "0000000000",
                                2512 => "0000001000",
                                2513 => "0000010000",
                                2514 => "0000010100",
                                2515 => "1011010000",
                                2516 => "1001110000",
                                2517 => "1011011000",
                                2518 => "1101000000",
                                2519 => "0001011100",
                                2520 => "0100101100",
                                2521 => "0000100100",
                                2522 => "0110000000",
                                2523 => "0011001000",
                                2524 => "1011000100",
                                2525 => "1000110000",
                                2526 => "0100011100",
                                2527 => "0100111100",
                                2528 => "0000100000",
                                2529 => "0000000000",
                                2530 => "0100010101",
                                2531 => "0100010110",
                                2532 => "0000000000",
                                2533 => "0000000000",
                                2534 => "0011000000",
                                2535 => "1100111000",
                                2536 => "1011100000",
                                2537 => "0100000000",
                                2538 => "0000000000",
                                2539 => "0110110000",
                                2540 => "0000011000",
                                2541 => "1101011100",
                                2542 => "0111000000",
                                2543 => "0011010000",
                                2544 => "1000111000",
                                2545 => "0111001000",
                                2546 => "0000001000",
                                2547 => "1100000000",
                                2548 => "1010100000",
                                2549 => "0000000100",
                                2550 => "0110011000",
                                2551 => "0000000100",
                                2552 => "1011101100",
                                2553 => "1110010000",
                                2554 => "1110110000",
                                2555 => "1000010000",
                                2556 => "1101001000",
                                2557 => "0100000100",
                                2558 => "1100000100",
                                2559 => "0000000000",
                                2560 => "1001010100",
                                2561 => "1001000000",
                                2562 => "0110011100",
                                2563 => "0111000000",
                                2564 => "0001001000",
                                2565 => "1111101000",
                                2566 => "1111000000",
                                2567 => "1110000100",
                                2568 => "0101101100",
                                2569 => "0000000000",
                                2570 => "0000000000",
                                2571 => "0000001000",
                                2572 => "0000010000",
                                2573 => "0000010100",
                                2574 => "1010000000",
                                2575 => "0000000100",
                                2576 => "0000000100",
                                2577 => "0000010000",
                                2578 => "0000001000",
                                2579 => "1001110000",
                                2580 => "1011011000",
                                2581 => "1101000000",
                                2582 => "0001011100",
                                2583 => "0100101100",
                                2584 => "0000100100",
                                2585 => "0110000000",
                                2586 => "0011001000",
                                2587 => "1011000100",
                                2588 => "1000110000",
                                2589 => "0100011100",
                                2590 => "0100111100",
                                2591 => "0000100000",
                                2592 => "0000000000",
                                2593 => "0100010101",
                                2594 => "0100010110",
                                2595 => "0000000000",
                                2596 => "0000000000",
                                2597 => "0011000000",
                                2598 => "0000000000",
                                2599 => "0000000000",
                                2600 => "0100000000",
                                2601 => "0000000000",
                                2602 => "1110010000",
                                2603 => "0000011000",
                                2604 => "0011011100",
                                2605 => "0010110100",
                                2606 => "0011010000",
                                2607 => "0001000100",
                                2608 => "0110100100",
                                2609 => "0111101100",
                                2610 => "1100000000",
                                2611 => "1010100000",
                                2612 => "0000000100",
                                2613 => "0110011000",
                                2614 => "0000000100",
                                2615 => "1011101100",
                                2616 => "1110010000",
                                2617 => "1110110100",
                                2618 => "0000010000",
                                2619 => "0010111100",
                                2620 => "0011010000",
                                2621 => "1111010100",
                                2622 => "1101110000",
                                2623 => "1011100000",
                                2624 => "0000000000",
                                2625 => "0100100000",
                                2626 => "0111000000",
                                2627 => "0001001000",
                                2628 => "0110100100",
                                2629 => "0000001100",
                                2630 => "1011110100",
                                2631 => "1010001100",
                                2632 => "0000000000",
                                2633 => "0000000000",
                                2634 => "0000001000",
                                2635 => "0000010000",
                                2636 => "0000010100",
                                2637 => "1011010000",
                                2638 => "0000000100",
                                2639 => "0000000100",
                                2640 => "0000010000",
                                2641 => "0000001000",
                                2642 => "1001110000",
                                2643 => "1011011000",
                                2644 => "1101000000",
                                2645 => "0001011100",
                                2646 => "0100101100",
                                2647 => "0000100100",
                                2648 => "0110000000",
                                2649 => "0011001000",
                                2650 => "1011000100",
                                2651 => "1000110000",
                                2652 => "0100011100",
                                2653 => "0100111100",
                                2654 => "0000100000",
                                2655 => "0000000000",
                                2656 => "0100010101",
                                2657 => "0100010110",
                                2658 => "0000000000",
                                2659 => "0000000000",
                                2660 => "0011000000",
                                2661 => "0100011100",
                                2662 => "0101000000",
                                2663 => "0100000000",
                                2664 => "0000000000",
                                2665 => "0110101000",
                                2666 => "0000011000",
                                2667 => "0011000000",
                                2668 => "1101101100",
                                2669 => "0010100000",
                                2670 => "0100110000",
                                2671 => "1010111000",
                                2672 => "0100001000",
                                2673 => "1100000000",
                                2674 => "1010100000",
                                2675 => "0000000100",
                                2676 => "0110011000",
                                2677 => "0000000100",
                                2678 => "1011101100",
                                2679 => "1110010000",
                                2680 => "1110101100",
                                2681 => "0001011100",
                                2682 => "1011100000",
                                2683 => "1011010100",
                                2684 => "1110100000",
                                2685 => "1110110100",
                                2686 => "0100010100",
                                2687 => "0010110000",
                                2688 => "0011001000",
                                2689 => "0111000000",
                                2690 => "0001001000",
                                2691 => "0010000000",
                                2692 => "0000000000",
                                2693 => "1111110000",
                                2694 => "1100011000",
                                2695 => "0000000000",
                                2696 => "0000000000",
                                2697 => "0000001000",
                                2698 => "0000010000",
                                2699 => "0000010100",
                                2700 => "1010000000",
                                2701 => "0000000100",
                                2702 => "0000000100",
                                2703 => "0000010000",
                                2704 => "0000001000",
                                2705 => "1001110000",
                                2706 => "1011011000",
                                2707 => "1101000000",
                                2708 => "0001011100",
                                2709 => "0100101100",
                                2710 => "0000100100",
                                2711 => "0110000000",
                                2712 => "0011001000",
                                2713 => "1011000100",
                                2714 => "1000110000",
                                2715 => "0100011100",
                                2716 => "0100111100",
                                2717 => "0000100000",
                                2718 => "0000000000",
                                2719 => "0100010101",
                                2720 => "0100010110",
                                2721 => "0000000000",
                                2722 => "0000000000",
                                2723 => "0011000000",
                                2724 => "0000000000",
                                2725 => "0000000000",
                                2726 => "0100000000",
                                2727 => "0000000000",
                                2728 => "0011100100",
                                2729 => "0000011000",
                                2730 => "1000110000",
                                2731 => "1111100000",
                                2732 => "1100011100",
                                2733 => "1110100000",
                                2734 => "0010101000",
                                2735 => "1101100100",
                                2736 => "1100000000",
                                2737 => "1010100000",
                                2738 => "0000000100",
                                2739 => "0110011000",
                                2740 => "0000000100",
                                2741 => "1011101100",
                                2742 => "1110010000",
                                2743 => "1110111000",
                                2744 => "1001101100",
                                2745 => "0100100100",
                                2746 => "0010111100",
                                2747 => "1010011000",
                                2748 => "1000010000",
                                2749 => "0000011100",
                                2750 => "0001111000",
                                2751 => "1000000100",
                                2752 => "0111000000",
                                2753 => "0001001000",
                                2754 => "1111111100",
                                2755 => "1111111100",
                                2756 => "0111101000",
                                2757 => "0001110100",
                                2758 => "0000000000",
                                2759 => "0000000000",
                                2760 => "0000001000",
                                2761 => "0000010000",
                                2762 => "0000010100",
                                2763 => "1011010000",
                                2764 => "0000000100",
                                2765 => "0000000100",
                                2766 => "0000010000",
                                2767 => "0000001000",
                                2768 => "1001110000",
                                2769 => "1011011000",
                                2770 => "1101000000",
                                2771 => "0001011100",
                                2772 => "0100101100",
                                2773 => "0000100100",
                                2774 => "0110000000",
                                2775 => "0011001000",
                                2776 => "1011000100",
                                2777 => "1000110000",
                                2778 => "0100011100",
                                2779 => "0100111100",
                                2780 => "0000100000",
                                2781 => "0000000000",
                                2782 => "0100010101",
                                2783 => "0100010110",
                                2784 => "0000000000",
                                2785 => "0000000000",
                                2786 => "0011000000",
                                2787 => "0001000100",
                                2788 => "0111010000",
                                2789 => "0000000000",
                                2790 => "0000000000",
                                2791 => "0011100000",
                                2792 => "0000011000",
                                2793 => "0100010000",
                                2794 => "0001101100",
                                2795 => "0000100000",
                                2796 => "1111110100",
                                2797 => "0110001000",
                                2798 => "0010111000",
                                2799 => "1100000000",
                                2800 => "1010100000",
                                2801 => "0000000100",
                                2802 => "0110011000",
                                2803 => "0000000100",
                                2804 => "1011101100",
                                2805 => "1110010000",
                                2806 => "1111000000",
                                2807 => "1011110000",
                                2808 => "1000101000",
                                2809 => "1011010100",
                                2810 => "0110000000",
                                2811 => "0000011000",
                                2812 => "1000110000",
                                2813 => "1101011100",
                                2814 => "0010111100",
                                2815 => "0111000000",
                                2816 => "0001001000",
                                2817 => "1111101000",
                                2818 => "1111000000",
                                2819 => "0010010000",
                                2820 => "1001001000",
                                2821 => "0000000000",
                                2822 => "0000000000",
                                2823 => "0000001000",
                                2824 => "0000010000",
                                2825 => "0000010100",
                                2826 => "1011010000",
                                2827 => "0000000100",
                                2828 => "0000000100",
                                2829 => "0000010000",
                                2830 => "0000001000",
                                2831 => "1001110000",
                                2832 => "1011011000",
                                2833 => "1101000000",
                                2834 => "0001011100",
                                2835 => "0100101100",
                                2836 => "0000100100",
                                2837 => "0110000000",
                                2838 => "0011001000",
                                2839 => "1011000100",
                                2840 => "1000110000",
                                2841 => "0100011100",
                                2842 => "0100111100",
                                2843 => "0000100000",
                                2844 => "0000000000",
                                2845 => "0100010101",
                                2846 => "0100010110",
                                2847 => "0000000000",
                                2848 => "0000000000",
                                2849 => "0011000000",
                                2850 => "0000000000",
                                2851 => "0000000000",
                                2852 => "0100000000",
                                2853 => "0000000000",
                                2854 => "0011010000",
                                2855 => "0000011000",
                                2856 => "1110001000",
                                2857 => "1000000000",
                                2858 => "1000100000",
                                2859 => "1111001100",
                                2860 => "0001100100",
                                2861 => "0100011000",
                                2862 => "1100000000",
                                2863 => "1010100000",
                                2864 => "0000000100",
                                2865 => "0110011000",
                                2866 => "0000000100",
                                2867 => "1011101100",
                                2868 => "1110010000",
                                2869 => "1110111100",
                                2870 => "0010010000",
                                2871 => "1110111000",
                                2872 => "0101101100",
                                2873 => "1100110000",
                                2874 => "1101111100",
                                2875 => "0001110100",
                                2876 => "1011001100",
                                2877 => "1100010000",
                                2878 => "0111000000",
                                2879 => "0001001000",
                                2880 => "1010010100",
                                2881 => "0110010000",
                                2882 => "0111111100",
                                2883 => "0001101100",
                                2884 => "0000000000",
                                2885 => "0000000000",
                                2886 => "0000001000",
                                2887 => "0000010000",
                                2888 => "0000010100",
                                2889 => "1011010000",
                                2890 => "0000000100",
                                2891 => "0000000100",
                                2892 => "0000010000",
                                2893 => "0000001000",
                                2894 => "1001110000",
                                2895 => "1011011000",
                                2896 => "1101000000",
                                2897 => "0001011100",
                                2898 => "0100101100",
                                2899 => "0000100100",
                                2900 => "0110000000",
                                2901 => "0011001000",
                                2902 => "1011000100",
                                2903 => "1000110000",
                                2904 => "0100011100",
                                2905 => "0100111100",
                                2906 => "0000100000",
                                2907 => "0000000000",
                                2908 => "0100010101",
                                2909 => "0100010110",
                                2910 => "0000000000",
                                2911 => "0000000000",
                                2912 => "0011000000",
                                2913 => "0100110000",
                                2914 => "1101100000",
                                2915 => "0000000000",
                                2916 => "0000000000",
                                2917 => "1111010000",
                                2918 => "0000011000",
                                2919 => "0011001100",
                                2920 => "1001111100",
                                2921 => "1000111100",
                                2922 => "1100110000",
                                2923 => "1111010000",
                                2924 => "0111010100",
                                2925 => "1100000000",
                                2926 => "1010100000",
                                2927 => "0000000100",
                                2928 => "0110011000",
                                2929 => "0000000100",
                                2930 => "1011101100",
                                2931 => "1110010000",
                                2932 => "1111000100",
                                2933 => "0000100100",
                                2934 => "1111001100",
                                2935 => "0000100000",
                                2936 => "1100110000",
                                2937 => "1000001000",
                                2938 => "0100100000",
                                2939 => "1101010000",
                                2940 => "0000110100",
                                2941 => "0111000000",
                                2942 => "0001001000",
                                2943 => "0000010100",
                                2944 => "1010000000",
                                2945 => "1110011100",
                                2946 => "0111000000",
                                2947 => "0000000000",
                                2948 => "0000000000",
                                2949 => "0000001000",
                                2950 => "0000010000",
                                2951 => "0000010100",
                                2952 => "1010000000",
                                2953 => "0000000100",
                                2954 => "0000000100",
                                2955 => "0000010000",
                                2956 => "0000001000",
                                2957 => "1001110000",
                                2958 => "1011011000",
                                2959 => "1101000000",
                                2960 => "0001011100",
                                2961 => "0100101100",
                                2962 => "0000100100",
                                2963 => "0110000000",
                                2964 => "0011001000",
                                2965 => "1011000100",
                                2966 => "1000110000",
                                2967 => "0100011100",
                                2968 => "0100111100",
                                2969 => "0000100000",
                                2970 => "0000000000",
                                2971 => "0100010101",
                                2972 => "0100010110",
                                2973 => "0000000000",
                                2974 => "0000000000",
                                2975 => "0011000000",
                                2976 => "1010001100",
                                2977 => "1011010000",
                                2978 => "0000000000",
                                2979 => "0000000000",
                                2980 => "1111001100",
                                2981 => "0000011000",
                                2982 => "1011110000",
                                2983 => "1000011100",
                                2984 => "0000110100",
                                2985 => "0010000100",
                                2986 => "1001100000",
                                2987 => "0101110000",
                                2988 => "1100000000",
                                2989 => "1010100000",
                                2990 => "0000000100",
                                2991 => "0110011000",
                                2992 => "0000000100",
                                2993 => "1011101100",
                                2994 => "1110010000",
                                2995 => "1111001000",
                                2996 => "0000111000",
                                2997 => "0110111000",
                                2998 => "0111111000",
                                2999 => "1000010000",
                                3000 => "1000011000",
                                3001 => "0111110000",
                                3002 => "1011011000",
                                3003 => "1000110000",
                                3004 => "0111000000",
                                3005 => "0001001000",
                                3006 => "0000010100",
                                3007 => "1010000000",
                                3008 => "0110010100",
                                3009 => "0100111000",
                                3010 => "0000000000",
                                3011 => "0000000000",
                                3012 => "0000001000",
                                3013 => "0000010000",
                                3014 => "0000010100",
                                3015 => "1010000000",
                                3016 => "0000000100",
                                3017 => "0000000100",
                                3018 => "0000010000",
                                3019 => "0000001000",
                                3020 => "1001110000",
                                3021 => "1011011000",
                                3022 => "1101000000",
                                3023 => "0001011100",
                                3024 => "0100101100",
                                3025 => "0000100100",
                                3026 => "0110000000",
                                3027 => "0011001000",
                                3028 => "1011000100",
                                3029 => "1000110000",
                                3030 => "0100011100",
                                3031 => "0100111100",
                                3032 => "0000100000",
                                3033 => "0000000000",
                                3034 => "0100010101",
                                3035 => "0100010110",
                                3036 => "0000000000",
                                3037 => "0000000000",
                                3038 => "0011000000",
                                3039 => "0000000000",
                                3040 => "0000000000",
                                3041 => "0100000000",
                                3042 => "0000000000",
                                3043 => "0011100000",
                                3044 => "0000011000",
                                3045 => "0110100100",
                                3046 => "0010001100",
                                3047 => "1001011100",
                                3048 => "1000101100",
                                3049 => "1000000000",
                                3050 => "0000101100",
                                3051 => "1100000000",
                                3052 => "1010100000",
                                3053 => "0000000100",
                                3054 => "0110011000",
                                3055 => "0000000100",
                                3056 => "1011101100",
                                3057 => "1110010000",
                                3058 => "1111001100",
                                3059 => "0000101100",
                                3060 => "0110001000",
                                3061 => "1111000100",
                                3062 => "0110010100",
                                3063 => "1111111100",
                                3064 => "0000111000",
                                3065 => "1110111000",
                                3066 => "0101110000",
                                3067 => "0111000000",
                                3068 => "0001001000",
                                3069 => "1111101000",
                                3070 => "1111000000",
                                3071 => "1101110100",
                                3072 => "1001011000",
                                3073 => "0000000000",
                                3074 => "0000000000",
                                3075 => "0000001000",
                                3076 => "0000010000",
                                3077 => "0000010100",
                                3078 => "1011010000",
                                3079 => "0000000100",
                                3080 => "0000000100",
                                3081 => "0000010000",
                                3082 => "0000001000",
                                3083 => "1001110000",
                                3084 => "1011011000",
                                3085 => "1101000000",
                                3086 => "0001011100",
                                3087 => "0100101100",
                                3088 => "0000100100",
                                3089 => "0110000000",
                                3090 => "0011001000",
                                3091 => "1011000100",
                                3092 => "1000110000",
                                3093 => "0100011100",
                                3094 => "0100111100",
                                3095 => "0000100000",
                                3096 => "0000000000",
                                3097 => "0100010101",
                                3098 => "0100010110",
                                3099 => "0000000000",
                                3100 => "0000000000",
                                3101 => "0011000000",
                                3102 => "0000101000",
                                3103 => "1000010100",
                                3104 => "0000000000",
                                3105 => "0000000000",
                                3106 => "0011100000",
                                3107 => "0000011000",
                                3108 => "0100101100",
                                3109 => "0000100000",
                                3110 => "0000100000",
                                3111 => "1111110100",
                                3112 => "0110001000",
                                3113 => "0011000000",
                                3114 => "1100000000",
                                3115 => "1010100000",
                                3116 => "0000000100",
                                3117 => "0110011000",
                                3118 => "0000000100",
                                3119 => "1011101100",
                                3120 => "1110010000",
                                3121 => "1111010000",
                                3122 => "1001010000",
                                3123 => "0001111000",
                                3124 => "0111110000",
                                3125 => "0110001000",
                                3126 => "0101010100",
                                3127 => "0110010100",
                                3128 => "1011110000",
                                3129 => "0001100100",
                                3130 => "0111000000",
                                3131 => "0001001000",
                                3132 => "1111101000",
                                3133 => "1111000000",
                                3134 => "0101001000",
                                3135 => "0011001100",
                                3136 => "0000000000",
                                3137 => "0000000000",
                                3138 => "0000001000",
                                3139 => "0000010000",
                                3140 => "0000010100",
                                3141 => "1011010000",
                                3142 => "0000000100",
                                3143 => "0000000100",
                                3144 => "0000010000",
                                3145 => "0000001000",
                                3146 => "1001110000",
                                3147 => "1011011000",
                                3148 => "1101000000",
                                3149 => "0001011100",
                                3150 => "0100101100",
                                3151 => "0000100100",
                                3152 => "0110000000",
                                3153 => "0011001000",
                                3154 => "1011000100",
                                3155 => "1000110000",
                                3156 => "0100011100",
                                3157 => "0100111100",
                                3158 => "0000100000",
                                3159 => "0000000000",
                                3160 => "0100010101",
                                3161 => "0100010110",
                                3162 => "0000000000",
                                3163 => "0000000000",
                                3164 => "0011000000",
                                3165 => "0001001100",
                                3166 => "0000001000",
                                3167 => "0000000000",
                                3168 => "0000000000",
                                3169 => "0011100000",
                                3170 => "0000011000",
                                3171 => "0100001000",
                                3172 => "1000110100",
                                3173 => "0000100000",
                                3174 => "1111110100",
                                3175 => "0110001000",
                                3176 => "0010111000",
                                3177 => "1100000000",
                                3178 => "1010100000",
                                3179 => "0000000100",
                                3180 => "0110011000",
                                3181 => "0000000100",
                                3182 => "1011101100",
                                3183 => "1110010000",
                                3184 => "1111010100",
                                3185 => "0001010100",
                                3186 => "1101010000",
                                3187 => "1110111100",
                                3188 => "0110100100",
                                3189 => "0000000000",
                                3190 => "1111111100",
                                3191 => "1100000000",
                                3192 => "1110001000",
                                3193 => "0111000000",
                                3194 => "0001001000",
                                3195 => "1111101000",
                                3196 => "1111000000",
                                3197 => "1010110100",
                                3198 => "0001010000",
                                3199 => "0000000000",
                                3200 => "0000000000",
                                3201 => "0000001000",
                                3202 => "0000010000",
                                3203 => "0000010100",
                                3204 => "1011010000",
                                3205 => "0000000100",
                                3206 => "0000000100",
                                3207 => "0000010000",
                                3208 => "0000001000",
                                3209 => "1001110000",
                                3210 => "1011011000",
                                3211 => "1101000000",
                                3212 => "0001011100",
                                3213 => "0100101100",
                                3214 => "0000100100",
                                3215 => "0110000000",
                                3216 => "0011001000",
                                3217 => "1011000100",
                                3218 => "1000110000",
                                3219 => "0100011100",
                                3220 => "0100111100",
                                3221 => "0000100000",
                                3222 => "0000000000",
                                3223 => "0100010101",
                                3224 => "0100010110",
                                3225 => "0000000000",
                                3226 => "0000000000",
                                3227 => "0011000000",
                                3228 => "1111101000",
                                3229 => "1001011100",
                                3230 => "0000000000",
                                3231 => "0000000000",
                                3232 => "0011100000",
                                3233 => "0000011000",
                                3234 => "0100111100",
                                3235 => "1011011100",
                                3236 => "0000100000",
                                3237 => "1111000100",
                                3238 => "0110110100",
                                3239 => "0111101000",
                                3240 => "1100000000",
                                3241 => "1010100000",
                                3242 => "0000000100",
                                3243 => "0110011000",
                                3244 => "0000000100",
                                3245 => "1011101100",
                                3246 => "1110010000",
                                3247 => "1111011000",
                                3248 => "1010000100",
                                3249 => "1111011100",
                                3250 => "0100001100",
                                3251 => "0100111100",
                                3252 => "0100101100",
                                3253 => "0110010000",
                                3254 => "1101011100",
                                3255 => "0110001100",
                                3256 => "0111000000",
                                3257 => "0001001000",
                                3258 => "1111101000",
                                3259 => "1111000000",
                                3260 => "0110000000",
                                3261 => "1110010000",
                                3262 => "0000000000",
                                3263 => "0000000000",
                                3264 => "0000001000",
                                3265 => "0000010000",
                                3266 => "0000010100",
                                3267 => "1011010000",
                                3268 => "0000000100",
                                3269 => "0000000100",
                                3270 => "0000010000",
                                3271 => "0000001000",
                                3272 => "1001110000",
                                3273 => "1011011000",
                                3274 => "1101000000",
                                3275 => "0001011100",
                                3276 => "0100101100",
                                3277 => "0000100100",
                                3278 => "0110000000",
                                3279 => "0011001000",
                                3280 => "1011000100",
                                3281 => "1000110000",
                                3282 => "0100011100",
                                3283 => "0100111100",
                                3284 => "0000100000",
                                3285 => "0000000000",
                                3286 => "0100010101",
                                3287 => "0100010110",
                                3288 => "0000000000",
                                3289 => "0000000000",
                                3290 => "0011000000",
                                3291 => "0000000000",
                                3292 => "0000000000",
                                3293 => "0100000000",
                                3294 => "0000000000",
                                3295 => "0011100000",
                                3296 => "0000011000",
                                3297 => "1000110100",
                                3298 => "1111100000",
                                3299 => "1100011100",
                                3300 => "1110100000",
                                3301 => "0010101000",
                                3302 => "1101100100",
                                3303 => "1100000000",
                                3304 => "1010100000",
                                3305 => "0000000100",
                                3306 => "0110011000",
                                3307 => "0000000100",
                                3308 => "1011101100",
                                3309 => "1110010000",
                                3310 => "1111011100",
                                3311 => "0000100100",
                                3312 => "1110110000",
                                3313 => "1000101100",
                                3314 => "1001100100",
                                3315 => "0110110100",
                                3316 => "1011001100",
                                3317 => "1000101100",
                                3318 => "0111110100",
                                3319 => "0111000000",
                                3320 => "0001001000",
                                3321 => "1111111100",
                                3322 => "1111111100",
                                3323 => "0101100000",
                                3324 => "1101011000",
                                3325 => "0000000000",
                                3326 => "0000000000",
                                3327 => "0000001000",
                                3328 => "0000010000",
                                3329 => "0000010100",
                                3330 => "1011010000",
                                3331 => "0000000100",
                                3332 => "0000000100",
                                3333 => "0000010000",
                                3334 => "0000001000",
                                3335 => "1001110000",
                                3336 => "1011011000",
                                3337 => "1101000000",
                                3338 => "0001011100",
                                3339 => "0100101100",
                                3340 => "0000100100",
                                3341 => "0110000000",
                                3342 => "0011001000",
                                3343 => "1011000100",
                                3344 => "1000110000",
                                3345 => "0100011100",
                                3346 => "0100111100",
                                3347 => "0000100000",
                                3348 => "0000000000",
                                3349 => "0100010101",
                                3350 => "0100010110",
                                3351 => "0000000000",
                                3352 => "0000000000",
                                3353 => "0010110000",
                                3354 => "0000000000",
                                3355 => "0000000000",
                                3356 => "0100000000",
                                3357 => "0000000000",
                                3358 => "1110010100",
                                3359 => "0000011000",
                                3360 => "1010110000",
                                3361 => "1000100100",
                                3362 => "0011011000",
                                3363 => "1110010100",
                                3364 => "1111000000",
                                3365 => "0100111000",
                                3366 => "1100000000",
                                3367 => "1010100000",
                                3368 => "0000000100",
                                3369 => "0110011000",
                                3370 => "0000000100",
                                3371 => "1011101100",
                                3372 => "1110010000",
                                3373 => "1111100000",
                                3374 => "1000000000",
                                3375 => "1101010000",
                                3376 => "1011001100",
                                3377 => "0000111000",
                                3378 => "0101100000",
                                3379 => "1000110000",
                                3380 => "1100100000",
                                3381 => "1011000000",
                                3382 => "0110000000",
                                3383 => "0001001000",
                                3384 => "0110100100",
                                3385 => "0000001100",
                                3386 => "0000100100",
                                3387 => "1111110100",
                                3388 => "0000000000",
                                3389 => "0000000000",
                                3390 => "0000001000",
                                3391 => "0000010000",
                                3392 => "0000010100",
                                3393 => "1011010000",
                                3394 => "1001110000",
                                3395 => "1011011000",
                                3396 => "1101000000",
                                3397 => "0001011100",
                                3398 => "0100101100",
                                3399 => "0000100100",
                                3400 => "0110000000",
                                3401 => "0011001000",
                                3402 => "1011000100",
                                3403 => "1000110000",
                                3404 => "0100011100",
                                3405 => "0100111100",
                                3406 => "0000100000",
                                3407 => "0000000000",
                                3408 => "0100010101",
                                3409 => "0100010110",
                                3410 => "0000000000",
                                3411 => "0000000000",
                                3412 => "0011000000",
                                3413 => "0000000000",
                                3414 => "0000000000",
                                3415 => "0100000000",
                                3416 => "0000000000",
                                3417 => "0011100000",
                                3418 => "0000011000",
                                3419 => "1000111000",
                                3420 => "1010000000",
                                3421 => "1100011100",
                                3422 => "1110100000",
                                3423 => "0010101000",
                                3424 => "0011000100",
                                3425 => "1100000000",
                                3426 => "1010100000",
                                3427 => "0000000100",
                                3428 => "0110011000",
                                3429 => "0000000100",
                                3430 => "1011101100",
                                3431 => "1110010000",
                                3432 => "1111100100",
                                3433 => "0000110000",
                                3434 => "0010001100",
                                3435 => "1011111000",
                                3436 => "0010000000",
                                3437 => "1101011100",
                                3438 => "0101010000",
                                3439 => "0101001000",
                                3440 => "1001011000",
                                3441 => "0111000000",
                                3442 => "0001001000",
                                3443 => "1111111100",
                                3444 => "1111111100",
                                3445 => "1111010000",
                                3446 => "0000001100",
                                3447 => "0000000000",
                                3448 => "0000000000",
                                3449 => "0000001000",
                                3450 => "0000010000",
                                3451 => "0000010100",
                                3452 => "1011010000",
                                3453 => "0000000100",
                                3454 => "0000000100",
                                3455 => "0000010000",
                                3456 => "0000001000",
                                3457 => "1001110000",
                                3458 => "1011011000",
                                3459 => "1101000000",
                                3460 => "0001011100",
                                3461 => "0100101100",
                                3462 => "0000100100",
                                3463 => "0110000000",
                                3464 => "0011001000",
                                3465 => "1011000100",
                                3466 => "1000110000",
                                3467 => "0100011100",
                                3468 => "0100111100",
                                3469 => "0000100000",
                                3470 => "0000000000",
                                3471 => "0100010101",
                                3472 => "0100010110",
                                3473 => "0000000000",
                                3474 => "0000000000",
                                3475 => "0011000000",
                                3476 => "0000000000",
                                3477 => "0000000000",
                                3478 => "0100000000",
                                3479 => "0000000000",
                                3480 => "0011001100",
                                3481 => "0000011000",
                                3482 => "0000111100",
                                3483 => "0001001000",
                                3484 => "0110100000",
                                3485 => "0001101000",
                                3486 => "0000111000",
                                3487 => "1000111000",
                                3488 => "1100000000",
                                3489 => "1010100000",
                                3490 => "0000000100",
                                3491 => "0110011000",
                                3492 => "0000000100",
                                3493 => "1011101100",
                                3494 => "1110010000",
                                3495 => "1111101000",
                                3496 => "1111010000",
                                3497 => "1101101100",
                                3498 => "1001001000",
                                3499 => "1011010000",
                                3500 => "0111011000",
                                3501 => "0001111000",
                                3502 => "0000001100",
                                3503 => "1001001000",
                                3504 => "0111000000",
                                3505 => "0001001000",
                                3506 => "1111111100",
                                3507 => "1111111100",
                                3508 => "0110001000",
                                3509 => "1001111000",
                                3510 => "0000000000",
                                3511 => "0000000000",
                                3512 => "0000001000",
                                3513 => "0000010000",
                                3514 => "0000010100",
                                3515 => "0111100000",
                                3516 => "0000000100",
                                3517 => "0000000100",
                                3518 => "0000010000",
                                3519 => "0000001000",
                                3520 => "1001110000",
                                3521 => "1011011000",
                                3522 => "1101000000",
                                3523 => "0001011100",
                                3524 => "0100101100",
                                3525 => "0000100100",
                                3526 => "0110000000",
                                3527 => "0011001000",
                                3528 => "1011000100",
                                3529 => "1000110000",
                                3530 => "0100011100",
                                3531 => "0100111100",
                                3532 => "0000100000",
                                3533 => "0000000000",
                                3534 => "0100010101",
                                3535 => "0100010110",
                                3536 => "0000000000",
                                3537 => "0000000000",
                                3538 => "0011000000",
                                3539 => "1000001100",
                                3540 => "0000000100",
                                3541 => "0000000000",
                                3542 => "0000000000",
                                3543 => "1111010000",
                                3544 => "0000011000",
                                3545 => "1111110100",
                                3546 => "1001111000",
                                3547 => "1000111100",
                                3548 => "1100110000",
                                3549 => "1111010000",
                                3550 => "0100110000",
                                3551 => "1100000000",
                                3552 => "1010100000",
                                3553 => "0000000100",
                                3554 => "0110011000",
                                3555 => "0000000100",
                                3556 => "1011101100",
                                3557 => "1110010000",
                                3558 => "1111101100",
                                3559 => "0000101000",
                                3560 => "0100000100",
                                3561 => "0001010000",
                                3562 => "0111000100",
                                3563 => "0000000100",
                                3564 => "0111001100",
                                3565 => "1011011100",
                                3566 => "0111101100",
                                3567 => "0111000000",
                                3568 => "0001001000",
                                3569 => "0000010100",
                                3570 => "1010000000",
                                3571 => "0111100100",
                                3572 => "0000010000",
                                3573 => "0000000000",
                                3574 => "0000000000",
                                3575 => "0000001000",
                                3576 => "0000010000",
                                3577 => "0000010100",
                                3578 => "1010000000",
                                3579 => "0000000100",
                                3580 => "0000000100",
                                3581 => "0000010000",
                                3582 => "0000001000",
                                3583 => "1001110000",
                                3584 => "1011011000",
                                3585 => "1101000000",
                                3586 => "0001011100",
                                3587 => "0100101100",
                                3588 => "0000100100",
                                3589 => "0110000000",
                                3590 => "0011001000",
                                3591 => "1011000100",
                                3592 => "1000110000",
                                3593 => "0100011100",
                                3594 => "0100111100",
                                3595 => "0000100000",
                                3596 => "0000000000",
                                3597 => "0100010101",
                                3598 => "0100010110",
                                3599 => "0000000000",
                                3600 => "0000000000",
                                3601 => "0011000000",
                                3602 => "0000000000",
                                3603 => "0000000000",
                                3604 => "0100000000",
                                3605 => "0000000000",
                                3606 => "0010100100",
                                3607 => "0000011000",
                                3608 => "0010000000",
                                3609 => "0001100100",
                                3610 => "0000111100",
                                3611 => "1011110000",
                                3612 => "0101111100",
                                3613 => "1110010100",
                                3614 => "1100000000",
                                3615 => "1010100000",
                                3616 => "0000000100",
                                3617 => "0110011000",
                                3618 => "0000000100",
                                3619 => "1011101100",
                                3620 => "1110010000",
                                3621 => "1111110000",
                                3622 => "0000111100",
                                3623 => "0110001000",
                                3624 => "0101101100",
                                3625 => "0001111000",
                                3626 => "0101010100",
                                3627 => "0110000000",
                                3628 => "0000110000",
                                3629 => "0100110100",
                                3630 => "0111000000",
                                3631 => "0001001000",
                                3632 => "1111111100",
                                3633 => "1111111100",
                                3634 => "1001111000",
                                3635 => "0111101000",
                                3636 => "0000000000",
                                3637 => "0000000000",
                                3638 => "0000001000",
                                3639 => "0000010000",
                                3640 => "0000010100",
                                3641 => "1011010000",
                                3642 => "0000000100",
                                3643 => "0000000100",
                                3644 => "0000010000",
                                3645 => "0000001000",
                                3646 => "1001110000",
                                3647 => "1011011000",
                                3648 => "1101000000",
                                3649 => "0001011100",
                                3650 => "0100101100",
                                3651 => "0000100100",
                                3652 => "0110000000",
                                3653 => "0011001000",
                                3654 => "1011000100",
                                3655 => "1000110000",
                                3656 => "0100011100",
                                3657 => "0100111100",
                                3658 => "0000100000",
                                3659 => "0000000000",
                                3660 => "0100010101",
                                3661 => "0100010110",
                                3662 => "0000000000",
                                3663 => "0000000000",
                                3664 => "0011000000",
                                3665 => "0000000000",
                                3666 => "0000000000",
                                3667 => "0100000000",
                                3668 => "0000000000",
                                3669 => "0011100000",
                                3670 => "0000011000",
                                3671 => "0101100000",
                                3672 => "0101100000",
                                3673 => "1011100100",
                                3674 => "1100011100",
                                3675 => "0110111000",
                                3676 => "1001101000",
                                3677 => "1100000000",
                                3678 => "1010100000",
                                3679 => "0000000100",
                                3680 => "0110011000",
                                3681 => "0000000100",
                                3682 => "1011101100",
                                3683 => "1110010000",
                                3684 => "1111110100",
                                3685 => "1100101100",
                                3686 => "1010100000",
                                3687 => "1010111000",
                                3688 => "0010100000",
                                3689 => "1001001000",
                                3690 => "0100010100",
                                3691 => "1011110100",
                                3692 => "0010011000",
                                3693 => "0111000000",
                                3694 => "0001001000",
                                3695 => "1111111100",
                                3696 => "1111111100",
                                3697 => "1110100000",
                                3698 => "1010100000",
                                3699 => "0000000000",
                                3700 => "0000000000",
                                3701 => "0000001000",
                                3702 => "0000010000",
                                3703 => "0000010100",
                                3704 => "1011010000",
                                3705 => "0000000100",
                                3706 => "0000000100",
                                3707 => "0000010000",
                                3708 => "0000001000",
                                3709 => "1001110000",
                                3710 => "1011011000",
                                3711 => "1101000000",
                                3712 => "0001011100",
                                3713 => "0100101100",
                                3714 => "0000100100",
                                3715 => "0110000000",
                                3716 => "0011001000",
                                3717 => "1011000100",
                                3718 => "1000110000",
                                3719 => "0100011100",
                                3720 => "0100111100",
                                3721 => "0000100000",
                                3722 => "0000000000",
                                3723 => "0100010101",
                                3724 => "0100010110",
                                3725 => "0000000000",
                                3726 => "0000000000",
                                3727 => "0011000000",
                                3728 => "0000000000",
                                3729 => "0000000000",
                                3730 => "0100000000",
                                3731 => "0000000000",
                                3732 => "0011001100",
                                3733 => "0000011000",
                                3734 => "1000000000",
                                3735 => "0110010000",
                                3736 => "1000110000",
                                3737 => "0101001000",
                                3738 => "0111100100",
                                3739 => "0000001100",
                                3740 => "1100000000",
                                3741 => "1010100000",
                                3742 => "0000000100",
                                3743 => "0110011000",
                                3744 => "0000000100",
                                3745 => "1011101100",
                                3746 => "1110010000",
                                3747 => "1111111000",
                                3748 => "1000000100",
                                3749 => "0100111100",
                                3750 => "1111100100",
                                3751 => "0010001100",
                                3752 => "1001111100",
                                3753 => "1100001100",
                                3754 => "0000110000",
                                3755 => "0010010100",
                                3756 => "0111000000",
                                3757 => "0001001000",
                                3758 => "1111111100",
                                3759 => "1111111100",
                                3760 => "1010111000",
                                3761 => "1010110100",
                                3762 => "0000000000",
                                3763 => "0000000000",
                                3764 => "0000001000",
                                3765 => "0000010000",
                                3766 => "0000010100",
                                3767 => "1001110000",
                                3768 => "0000000100",
                                3769 => "0000000100",
                                3770 => "0000010000",
                                3771 => "0000001000",
                                3772 => "1001110000",
                                3773 => "1011011000",
                                3774 => "1101000000",
                                3775 => "0001011100",
                                3776 => "0100101100",
                                3777 => "0000100100",
                                3778 => "0110000000",
                                3779 => "0011001000",
                                3780 => "1011000100",
                                3781 => "1000110000",
                                3782 => "0100011100",
                                3783 => "0100111100",
                                3784 => "0000100000",
                                3785 => "0000000000",
                                3786 => "0100010101",
                                3787 => "0100010110",
                                3788 => "0000000000",
                                3789 => "0000000000",
                                3790 => "0011000000",
                                3791 => "0000000000",
                                3792 => "0000000000",
                                3793 => "0100000000",
                                3794 => "0000000000",
                                3795 => "1111000000",
                                3796 => "0000011000",
                                3797 => "1100101100",
                                3798 => "0001010100",
                                3799 => "0010001100",
                                3800 => "1001110000",
                                3801 => "1101101000",
                                3802 => "0000011100",
                                3803 => "1100000000",
                                3804 => "1010100000",
                                3805 => "0000000100",
                                3806 => "0110011000",
                                3807 => "0000000100",
                                3808 => "1011101100",
                                3809 => "1110010000",
                                3810 => "1111111100",
                                3811 => "1101110000",
                                3812 => "1001000100",
                                3813 => "1111001100",
                                3814 => "0101110000",
                                3815 => "1000000100",
                                3816 => "1111010000",
                                3817 => "1110010000",
                                3818 => "1001000000",
                                3819 => "0111000000",
                                3820 => "0001001000",
                                3821 => "0110100100",
                                3822 => "0000001100",
                                3823 => "0011110100",
                                3824 => "0010101100",
                                3825 => "0000000000",
                                3826 => "0000000000",
                                3827 => "0000001000",
                                3828 => "0000010000",
                                3829 => "0000010100",
                                3830 => "1011010000",
                                3831 => "0000000100",
                                3832 => "0000000100",
                                3833 => "0000010000",
                                3834 => "0000001000",
                                3835 => "1001110000",
                                3836 => "1011011000",
                                3837 => "1101000000",
                                3838 => "0001011100",
                                3839 => "0100101100",
                                3840 => "0000100100",
                                3841 => "0110000000",
                                3842 => "0011001000",
                                3843 => "1011000100",
                                3844 => "1000110000",
                                3845 => "0100011100",
                                3846 => "0100111100",
                                3847 => "0000100000",
                                3848 => "0000000000",
                                3849 => "0100010101",
                                3850 => "0100010110",
                                3851 => "0000000000",
                                3852 => "0000000000",
                                3853 => "0011000000",
                                3854 => "0111010000",
                                3855 => "1100010100",
                                3856 => "0100000000",
                                3857 => "0000000000",
                                3858 => "1110100000",
                                3859 => "0000011000",
                                3860 => "0010110100",
                                3861 => "1110001000",
                                3862 => "1000111000",
                                3863 => "0000000000",
                                3864 => "1010000000",
                                3865 => "0001000100",
                                3866 => "1100000000",
                                3867 => "1010100000",
                                3868 => "0000000100",
                                3869 => "0110011000",
                                3870 => "0000000100",
                                3871 => "1011101100",
                                3872 => "1110010100",
                                3873 => "0000000000",
                                3874 => "1010000000",
                                3875 => "1000011000",
                                3876 => "0011101100",
                                3877 => "1111010000",
                                3878 => "1100011100",
                                3879 => "0100101100",
                                3880 => "1100111000",
                                3881 => "0011001100",
                                3882 => "0111000000",
                                3883 => "0001001000",
                                3884 => "0011010000",
                                3885 => "1011110000",
                                3886 => "0000011000",
                                3887 => "1110110000",
                                3888 => "0000000000",
                                3889 => "0000000000",
                                3890 => "0000001000",
                                3891 => "0000010000",
                                3892 => "0000010100",
                                3893 => "0100011000",
                                3894 => "0000010000",
                                3895 => "0000001000",
                                3896 => "0000000000",
                                3897 => "0000000000",
                                3898 => "1001110000",
                                3899 => "1011011000",
                                3900 => "1101000000",
                                3901 => "0001011100",
                                3902 => "0100101100",
                                3903 => "0000100100",
                                3904 => "0110000000",
                                3905 => "0011001000",
                                3906 => "1011000100",
                                3907 => "1000110000",
                                3908 => "0100011100",
                                3909 => "0100111100",
                                3910 => "0000100000",
                                3911 => "0000000000",
                                3912 => "0100010101",
                                3913 => "0100010110",
                                3914 => "0000000000",
                                3915 => "0000000000",
                                3916 => "0011000000",
                                3917 => "1111111000",
                                3918 => "0010010100",
                                3919 => "0100000000",
                                3920 => "0000000000",
                                3921 => "1110011100",
                                3922 => "0000011000",
                                3923 => "1010010100",
                                3924 => "1000000100",
                                3925 => "1000111000",
                                3926 => "0000000000",
                                3927 => "1010000000",
                                3928 => "0001000100",
                                3929 => "1100000000",
                                3930 => "1010100000",
                                3931 => "0000000100",
                                3932 => "0110011000",
                                3933 => "0000000100",
                                3934 => "1011101100",
                                3935 => "1110010100",
                                3936 => "0000000100",
                                3937 => "0111100100",
                                3938 => "0101000100",
                                3939 => "0110000000",
                                3940 => "0010010000",
                                3941 => "0001100100",
                                3942 => "0011011100",
                                3943 => "0110110000",
                                3944 => "0000010100",
                                3945 => "0111000000",
                                3946 => "0001001000",
                                3947 => "0011010000",
                                3948 => "1011110000",
                                3949 => "0001101000",
                                3950 => "0011001100",
                                3951 => "0000000000",
                                3952 => "0000000000",
                                3953 => "0000001000",
                                3954 => "0000010000",
                                3955 => "0000010100",
                                3956 => "0100011000",
                                3957 => "0000010000",
                                3958 => "0000001000",
                                3959 => "0000000000",
                                3960 => "0000000000",
                                3961 => "1001110000",
                                3962 => "1011011000",
                                3963 => "1101000000",
                                3964 => "0001011100",
                                3965 => "0100101100",
                                3966 => "0000100100",
                                3967 => "0110000000",
                                3968 => "0011001000",
                                3969 => "1011000100",
                                3970 => "1000110000",
                                3971 => "0100011100",
                                3972 => "0100111100",
                                3973 => "0000100000",
                                3974 => "0000000000",
                                3975 => "0100010101",
                                3976 => "0100010110",
                                3977 => "0000000000",
                                3978 => "0000000000",
                                3979 => "0011000000",
                                3980 => "0000000000",
                                3981 => "0000000000",
                                3982 => "0100000000",
                                3983 => "0000000000",
                                3984 => "1110010000",
                                3985 => "0000011000",
                                3986 => "0100011100",
                                3987 => "1110100000",
                                3988 => "0011010000",
                                3989 => "0011001100",
                                3990 => "0101100000",
                                3991 => "1001111000",
                                3992 => "1100000000",
                                3993 => "1010100000",
                                3994 => "0000000100",
                                3995 => "0110011000",
                                3996 => "0000000100",
                                3997 => "1011101100",
                                3998 => "1110010100",
                                3999 => "0000001000",
                                4000 => "1000110100",
                                4001 => "0110000100",
                                4002 => "1101010000",
                                4003 => "0011110000",
                                4004 => "1000111000",
                                4005 => "1110001100",
                                4006 => "1110010000",
                                4007 => "1000010000",
                                4008 => "0111000000",
                                4009 => "0001001000",
                                4010 => "0110100100",
                                4011 => "0000001100",
                                4012 => "0000111100",
                                4013 => "0110100000",
                                4014 => "0000000000",
                                4015 => "0000000000",
                                4016 => "0000001000",
                                4017 => "0000010000",
                                4018 => "0000010100",
                                4019 => "1011010000",
                                4020 => "0000000100",
                                4021 => "0000000100",
                                4022 => "0000010000",
                                4023 => "0000001000",
                                4024 => "1001110000",
                                4025 => "1011011000",
                                4026 => "1101000000",
                                4027 => "0001011100",
                                4028 => "0100101100",
                                4029 => "0000100100",
                                4030 => "0110000000",
                                4031 => "0011001000",
                                4032 => "1011000100",
                                4033 => "1000110000",
                                4034 => "0100011100",
                                4035 => "0100111100",
                                4036 => "0000100000",
                                4037 => "0000000000",
                                4038 => "0100010101",
                                4039 => "0100010110",
                                4040 => "0000000000",
                                4041 => "0000000000",
                                4042 => "0011000000",
                                4043 => "0000000000",
                                4044 => "0000000000",
                                4045 => "0100000000",
                                4046 => "0000000000",
                                4047 => "0010111100",
                                4048 => "0000011000",
                                4049 => "1010110000",
                                4050 => "1101100100",
                                4051 => "1000011000",
                                4052 => "1110000000",
                                4053 => "0101011000",
                                4054 => "0000000000",
                                4055 => "1100000000",
                                4056 => "1010100000",
                                4057 => "0000000100",
                                4058 => "0110011000",
                                4059 => "0000000100",
                                4060 => "1011101100",
                                4061 => "1110010100",
                                4062 => "0000010000",
                                4063 => "0000000100",
                                4064 => "1100100100",
                                4065 => "1111000100",
                                4066 => "0111110100",
                                4067 => "1100001000",
                                4068 => "1101100100",
                                4069 => "1011001000",
                                4070 => "1100110100",
                                4071 => "0111000000",
                                4072 => "0001001000",
                                4073 => "0110100100",
                                4074 => "0000001100",
                                4075 => "0010101100",
                                4076 => "0110111100",
                                4077 => "0000000000",
                                4078 => "0000000000",
                                4079 => "0000001000",
                                4080 => "0000010000",
                                4081 => "0000010100",
                                4082 => "1011010000",
                                4083 => "0000000100",
                                4084 => "0000000100",
                                4085 => "0000010000",
                                4086 => "0000001000",
                                4087 => "1001110000",
                                4088 => "1011011000",
                                4089 => "1101000000",
                                4090 => "0001011100",
                                4091 => "0100101100",
                                4092 => "0000100100",
                                4093 => "0110000000",
                                4094 => "0011001000",
                                4095 => "1011000100",
                                4096 => "1000110000",
                                4097 => "0100011100",
                                4098 => "0100111100",
                                4099 => "0000100000",
                                4100 => "0000000000",
                                4101 => "0100010101",
                                4102 => "0100010110",
                                4103 => "0000000000",
                                4104 => "0000000000",
                                4105 => "0011000000",
                                4106 => "0000000000",
                                4107 => "0000000000",
                                4108 => "0100000000",
                                4109 => "0000000000",
                                4110 => "1110010000",
                                4111 => "0000011000",
                                4112 => "1101111000",
                                4113 => "1110010000",
                                4114 => "0011010000",
                                4115 => "0001001000",
                                4116 => "1100000100",
                                4117 => "1100001000",
                                4118 => "1100000000",
                                4119 => "1010100000",
                                4120 => "0000000100",
                                4121 => "0110011000",
                                4122 => "0000000100",
                                4123 => "1011101100",
                                4124 => "1110010100",
                                4125 => "0000001100",
                                4126 => "0011010000",
                                4127 => "1111011100",
                                4128 => "0000010000",
                                4129 => "0111000100",
                                4130 => "0100111000",
                                4131 => "0111111000",
                                4132 => "0111101100",
                                4133 => "0100011100",
                                4134 => "0111000000",
                                4135 => "0001001000",
                                4136 => "0110100100",
                                4137 => "0000001100",
                                4138 => "0111100000",
                                4139 => "0011110000",
                                4140 => "0000000000",
                                4141 => "0000000000",
                                4142 => "0000001000",
                                4143 => "0000010000",
                                4144 => "0000010100",
                                4145 => "1011010000",
                                4146 => "0000000100",
                                4147 => "0000000100",
                                4148 => "0000010000",
                                4149 => "0000001000",
                                4150 => "1001110000",
                                4151 => "1011011000",
                                4152 => "1101000000",
                                4153 => "0001011100",
                                4154 => "0100101100",
                                4155 => "0000100100",
                                4156 => "0110000000",
                                4157 => "0011001000",
                                4158 => "1011000100",
                                4159 => "1000110000",
                                4160 => "0100011100",
                                4161 => "0100111100",
                                4162 => "0000100000",
                                4163 => "0000000000",
                                4164 => "0100010101",
                                4165 => "0100010110",
                                4166 => "0000000000",
                                4167 => "0000000000",
                                4168 => "0011000000",
                                4169 => "0000100000",
                                4170 => "1010011100",
                                4171 => "0000000000",
                                4172 => "0000000000",
                                4173 => "1111001100",
                                4174 => "0000011000",
                                4175 => "0101011100",
                                4176 => "1011101100",
                                4177 => "0000110100",
                                4178 => "0010000100",
                                4179 => "1001100000",
                                4180 => "0011011000",
                                4181 => "1100000000",
                                4182 => "1010100000",
                                4183 => "0000000100",
                                4184 => "0110011000",
                                4185 => "0000000100",
                                4186 => "1011101100",
                                4187 => "1110010100",
                                4188 => "0000010100",
                                4189 => "1010101100",
                                4190 => "0000011000",
                                4191 => "0000100100",
                                4192 => "1000000100",
                                4193 => "1010000000",
                                4194 => "1010111100",
                                4195 => "1101100100",
                                4196 => "0001001000",
                                4197 => "0111000000",
                                4198 => "0001001000",
                                4199 => "0000010100",
                                4200 => "1010000000",
                                4201 => "0000000100",
                                4202 => "0001001100",
                                4203 => "0000000000",
                                4204 => "0000000000",
                                4205 => "0000001000",
                                4206 => "0000010000",
                                4207 => "0000010100",
                                4208 => "1010000000",
                                4209 => "0000000100",
                                4210 => "0000000100",
                                4211 => "0000010000",
                                4212 => "0000001000",
                                4213 => "1001110000",
                                4214 => "1011011000",
                                4215 => "1101000000",
                                4216 => "0001011100",
                                4217 => "0100101100",
                                4218 => "0000100100",
                                4219 => "0110000000",
                                4220 => "0011001000",
                                4221 => "1011000100",
                                4222 => "1000110000",
                                4223 => "0100011100",
                                4224 => "0100111100",
                                4225 => "0000100000",
                                4226 => "0000000000",
                                4227 => "0100010101",
                                4228 => "0100010110",
                                4229 => "0000000000",
                                4230 => "0000000000",
                                4231 => "0011000000",
                                4232 => "0000000000",
                                4233 => "0000000000",
                                4234 => "0100000000",
                                4235 => "0000000000",
                                4236 => "0011100000",
                                4237 => "0000011000",
                                4238 => "1111110100",
                                4239 => "0100010100",
                                4240 => "0110100000",
                                4241 => "0101111000",
                                4242 => "0001101100",
                                4243 => "0001011000",
                                4244 => "1100000000",
                                4245 => "1010100000",
                                4246 => "0000000100",
                                4247 => "0110011000",
                                4248 => "0000000100",
                                4249 => "1011101100",
                                4250 => "1110010100",
                                4251 => "0000011000",
                                4252 => "0110010000",
                                4253 => "1110110100",
                                4254 => "0111000000",
                                4255 => "1011011100",
                                4256 => "1100001100",
                                4257 => "0100111000",
                                4258 => "0011100000",
                                4259 => "0111110100",
                                4260 => "0111000000",
                                4261 => "0001001000",
                                4262 => "1111101000",
                                4263 => "1111000000",
                                4264 => "1000101000",
                                4265 => "0110100100",
                                4266 => "0000000000",
                                4267 => "0000000000",
                                4268 => "0000001000",
                                4269 => "0000010000",
                                4270 => "0000010100",
                                4271 => "1011010000",
                                4272 => "0000000100",
                                4273 => "0000000100",
                                4274 => "0000010000",
                                4275 => "0000001000",
                                4276 => "1001110000",
                                4277 => "1011011000",
                                4278 => "1101000000",
                                4279 => "0001011100",
                                4280 => "0100101100",
                                4281 => "0000100100",
                                4282 => "0110000000",
                                4283 => "0011001000",
                                4284 => "1011000100",
                                4285 => "1000110000",
                                4286 => "0100011100",
                                4287 => "0100111100",
                                4288 => "0000100000",
                                4289 => "0000000000",
                                4290 => "0100010101",
                                4291 => "0100010110",
                                4292 => "0000000000",
                                4293 => "0000000000",
                                4294 => "0011000000",
                                4295 => "0000000000",
                                4296 => "0000000000",
                                4297 => "0100000000",
                                4298 => "0000000000",
                                4299 => "0011100100",
                                4300 => "0000011000",
                                4301 => "0101011100",
                                4302 => "0101100000",
                                4303 => "1011100100",
                                4304 => "1100011100",
                                4305 => "0110111000",
                                4306 => "1001101000",
                                4307 => "1100000000",
                                4308 => "1010100000",
                                4309 => "0000000100",
                                4310 => "0110011000",
                                4311 => "0000000100",
                                4312 => "1011101100",
                                4313 => "1110010100",
                                4314 => "0000011100",
                                4315 => "0100111100",
                                4316 => "1010000100",
                                4317 => "1011100000",
                                4318 => "0100111000",
                                4319 => "1011001000",
                                4320 => "1000001100",
                                4321 => "0111100000",
                                4322 => "1010111000",
                                4323 => "0111000000",
                                4324 => "0001001000",
                                4325 => "1111111100",
                                4326 => "1111111100",
                                4327 => "0111111000",
                                4328 => "1011101000",
                                4329 => "0000000000",
                                4330 => "0000000000",
                                4331 => "0000001000",
                                4332 => "0000010000",
                                4333 => "0000010100",
                                4334 => "1011010000",
                                4335 => "0000000100",
                                4336 => "0000000100",
                                4337 => "0000010000",
                                4338 => "0000001000",
                                4339 => "1001110000",
                                4340 => "1011011000",
                                4341 => "1101000000",
                                4342 => "0001011100",
                                4343 => "0100101100",
                                4344 => "0000100100",
                                4345 => "0110000000",
                                4346 => "0011001000",
                                4347 => "1011000100",
                                4348 => "1000110000",
                                4349 => "0100011100",
                                4350 => "0100111100",
                                4351 => "0000100000",
                                4352 => "0000000000",
                                4353 => "0100010101",
                                4354 => "0100010110",
                                4355 => "0000000000",
                                4356 => "0000000000",
                                4357 => "0011000000",
                                4358 => "0000000000",
                                4359 => "0000000000",
                                4360 => "0100000000",
                                4361 => "0000000000",
                                4362 => "0011100000",
                                4363 => "0000011000",
                                4364 => "0101101000",
                                4365 => "0110110100",
                                4366 => "1011100100",
                                4367 => "1100011100",
                                4368 => "0110110000",
                                4369 => "1000010100",
                                4370 => "1100000000",
                                4371 => "1010100000",
                                4372 => "0000000100",
                                4373 => "0110011000",
                                4374 => "0000000100",
                                4375 => "1011101100",
                                4376 => "1110010100",
                                4377 => "0000100000",
                                4378 => "0010101100",
                                4379 => "1000100000",
                                4380 => "1010000100",
                                4381 => "1110000100",
                                4382 => "0011110100",
                                4383 => "0000000100",
                                4384 => "0011000100",
                                4385 => "1100000100",
                                4386 => "0111000000",
                                4387 => "0001001000",
                                4388 => "1111111100",
                                4389 => "1111111100",
                                4390 => "0111011100",
                                4391 => "1100010000",
                                4392 => "0000000000",
                                4393 => "0000000000",
                                4394 => "0000001000",
                                4395 => "0000010000",
                                4396 => "0000010100",
                                4397 => "1011010000",
                                4398 => "0000000100",
                                4399 => "0000000100",
                                4400 => "0000010000",
                                4401 => "0000001000",
                                4402 => "1001110000",
                                4403 => "1011011000",
                                4404 => "1101000000",
                                4405 => "0001011100",
                                4406 => "0100101100",
                                4407 => "0000100100",
                                4408 => "0110000000",
                                4409 => "0011001000",
                                4410 => "1011000100",
                                4411 => "1000110000",
                                4412 => "0100011100",
                                4413 => "0100111100",
                                4414 => "0000100000",
                                4415 => "0000000000",
                                4416 => "0100010101",
                                4417 => "0100010110",
                                4418 => "0000000000",
                                4419 => "0000000000",
                                4420 => "0011000000",
                                4421 => "0000000000",
                                4422 => "0000000000",
                                4423 => "0100000000",
                                4424 => "0000000000",
                                4425 => "0011100100",
                                4426 => "0000011000",
                                4427 => "1000001100",
                                4428 => "0110100100",
                                4429 => "0110100000",
                                4430 => "0001000000",
                                4431 => "1001010000",
                                4432 => "0100000000",
                                4433 => "1100000000",
                                4434 => "1010100000",
                                4435 => "0000000100",
                                4436 => "0110011000",
                                4437 => "0000000100",
                                4438 => "1011101100",
                                4439 => "1110010100",
                                4440 => "0000100100",
                                4441 => "1001000100",
                                4442 => "1000101000",
                                4443 => "0010101100",
                                4444 => "1000010100",
                                4445 => "1101001000",
                                4446 => "0101001100",
                                4447 => "0100010000",
                                4448 => "1110100100",
                                4449 => "0111000000",
                                4450 => "0001001000",
                                4451 => "1111111100",
                                4452 => "1111111100",
                                4453 => "0000100100",
                                4454 => "1101101100",
                                4455 => "0000000000",
                                4456 => "0000000000",
                                4457 => "0000001000",
                                4458 => "0000010000",
                                4459 => "0000010100",
                                4460 => "0111100000",
                                4461 => "0000000100",
                                4462 => "0000000100",
                                4463 => "0000010000",
                                4464 => "0000001000",
                                4465 => "1001110000",
                                4466 => "1011011000",
                                4467 => "1101000000",
                                4468 => "0001011100",
                                4469 => "0100101100",
                                4470 => "0000100100",
                                4471 => "0110000000",
                                4472 => "0011001000",
                                4473 => "1011000100",
                                4474 => "1000110000",
                                4475 => "0100011100",
                                4476 => "0100111100",
                                4477 => "0000100000",
                                4478 => "0000000000",
                                4479 => "0100010101",
                                4480 => "0100010110",
                                4481 => "0000000000",
                                4482 => "0000000000",
                                4483 => "0011000000",
                                4484 => "0000000000",
                                4485 => "0000000000",
                                4486 => "0100000000",
                                4487 => "0000000000",
                                4488 => "0011100100",
                                4489 => "0000011000",
                                4490 => "1000001100",
                                4491 => "0110100100",
                                4492 => "0110100000",
                                4493 => "0001000000",
                                4494 => "1001010000",
                                4495 => "0100000000",
                                4496 => "1100000000",
                                4497 => "1010100000",
                                4498 => "0000000100",
                                4499 => "0110011000",
                                4500 => "0000000100",
                                4501 => "1011101100",
                                4502 => "1110010100",
                                4503 => "0000101000",
                                4504 => "0101010100",
                                4505 => "1000101000",
                                4506 => "0000111100",
                                4507 => "1010000000",
                                4508 => "1001001100",
                                4509 => "1001100000",
                                4510 => "0111011000",
                                4511 => "0111000100",
                                4512 => "0111000000",
                                4513 => "0001001000",
                                4514 => "1111111100",
                                4515 => "1111111100",
                                4516 => "0110111000",
                                4517 => "1111001000",
                                4518 => "0000000000",
                                4519 => "0000000000",
                                4520 => "0000001000",
                                4521 => "0000010000",
                                4522 => "0000010100",
                                4523 => "0111100000",
                                4524 => "0000000100",
                                4525 => "0000000100",
                                4526 => "0000010000",
                                4527 => "0000001000",
                                4528 => "1001110000",
                                4529 => "1011011000",
                                4530 => "1101000000",
                                4531 => "0001011100",
                                4532 => "0100101100",
                                4533 => "0000100100",
                                4534 => "0110000000",
                                4535 => "0011001000",
                                4536 => "1011000100",
                                4537 => "1000110000",
                                4538 => "0100011100",
                                4539 => "0100111100",
                                4540 => "0000100000",
                                4541 => "0000000000",
                                4542 => "0100010101",
                                4543 => "0100010110",
                                4544 => "0000000000",
                                4545 => "0000000000",
                                4546 => "0011000000",
                                4547 => "1110000100",
                                4548 => "1111010000",
                                4549 => "0000000000",
                                4550 => "0000000000",
                                4551 => "1111010000",
                                4552 => "0000011000",
                                4553 => "0111110100",
                                4554 => "0010111100",
                                4555 => "0000110100",
                                4556 => "0010000100",
                                4557 => "1001100000",
                                4558 => "0111010000",
                                4559 => "1100000000",
                                4560 => "1010100000",
                                4561 => "0000000100",
                                4562 => "0110011000",
                                4563 => "0000000100",
                                4564 => "1011101100",
                                4565 => "1110010100",
                                4566 => "0000101100",
                                4567 => "0001001000",
                                4568 => "1011010100",
                                4569 => "1000111000",
                                4570 => "0110111000",
                                4571 => "1111011100",
                                4572 => "0100000000",
                                4573 => "1000011100",
                                4574 => "1000011100",
                                4575 => "0111000000",
                                4576 => "0001001000",
                                4577 => "0000010100",
                                4578 => "1010000000",
                                4579 => "0000111100",
                                4580 => "0010110100",
                                4581 => "0000000000",
                                4582 => "0000000000",
                                4583 => "0000001000",
                                4584 => "0000010000",
                                4585 => "0000010100",
                                4586 => "1010000000",
                                4587 => "0000000100",
                                4588 => "0000000100",
                                4589 => "0000010000",
                                4590 => "0000001000",
                                4591 => "1001110000",
                                4592 => "1011011000",
                                4593 => "1101000000",
                                4594 => "0001011100",
                                4595 => "0100101100",
                                4596 => "0000100100",
                                4597 => "0110000000",
                                4598 => "0011001000",
                                4599 => "1011000100",
                                4600 => "1000110000",
                                4601 => "0100011100",
                                4602 => "0100111100",
                                4603 => "0000100000",
                                4604 => "0000000000",
                                4605 => "0100010101",
                                4606 => "0100010110",
                                4607 => "0000000000",
                                4608 => "0000000000",
                                4609 => "0011000000",
                                4610 => "1011101000",
                                4611 => "0101100100",
                                4612 => "0000000000",
                                4613 => "0000000000",
                                4614 => "1111001100",
                                4615 => "0000011000",
                                4616 => "1100011100",
                                4617 => "0100010100",
                                4618 => "1000111100",
                                4619 => "1100110000",
                                4620 => "1111010000",
                                4621 => "0100110100",
                                4622 => "1100000000",
                                4623 => "1010100000",
                                4624 => "0000000100",
                                4625 => "0110011000",
                                4626 => "0000000100",
                                4627 => "1011101100",
                                4628 => "1110010100",
                                4629 => "0000110000",
                                4630 => "1111100000",
                                4631 => "0100001100",
                                4632 => "1101111100",
                                4633 => "0100011100",
                                4634 => "1100100100",
                                4635 => "0000001100",
                                4636 => "0100111100",
                                4637 => "0000101000",
                                4638 => "0111000000",
                                4639 => "0001001000",
                                4640 => "0000010100",
                                4641 => "1010000000",
                                4642 => "0110000000",
                                4643 => "1111100100",
                                4644 => "0000000000",
                                4645 => "0000000000",
                                4646 => "0000001000",
                                4647 => "0000010000",
                                4648 => "0000010100",
                                4649 => "1010000000",
                                4650 => "0000000100",
                                4651 => "0000000100",
                                4652 => "0000010000",
                                4653 => "0000001000",
                                4654 => "1001110000",
                                4655 => "1011011000",
                                4656 => "1101000000",
                                4657 => "0001011100",
                                4658 => "0100101100",
                                4659 => "0000100100",
                                4660 => "0110000000",
                                4661 => "0011001000",
                                4662 => "1011000100",
                                4663 => "1000110000",
                                4664 => "0100011100",
                                4665 => "0100111100",
                                4666 => "0000100000",
                                4667 => "0000000000",
                                4668 => "0100010101",
                                4669 => "0100010110",
                                4670 => "0000000000",
                                4671 => "0000000000",
                                4672 => "0011000000",
                                4673 => "1011101000",
                                4674 => "0101101100",
                                4675 => "0000000000",
                                4676 => "0000000000",
                                4677 => "1111001100",
                                4678 => "0000011000",
                                4679 => "1100011100",
                                4680 => "0100001100",
                                4681 => "1000111100",
                                4682 => "1100110000",
                                4683 => "1111010000",
                                4684 => "0100110100",
                                4685 => "1100000000",
                                4686 => "1010100000",
                                4687 => "0000000100",
                                4688 => "0110011000",
                                4689 => "0000000100",
                                4690 => "1011101100",
                                4691 => "1110010100",
                                4692 => "0000110000",
                                4693 => "1111100000",
                                4694 => "0100001100",
                                4695 => "1101111100",
                                4696 => "0100011100",
                                4697 => "1100100100",
                                4698 => "0000001100",
                                4699 => "0100111100",
                                4700 => "0000101000",
                                4701 => "0111000000",
                                4702 => "0001001000",
                                4703 => "0000010100",
                                4704 => "1010000000",
                                4705 => "0110000000",
                                4706 => "1111100100",
                                4707 => "0000000000",
                                4708 => "0000000000",
                                4709 => "0000001000",
                                4710 => "0000010000",
                                4711 => "0000010100",
                                4712 => "1010000000",
                                4713 => "0000000100",
                                4714 => "0000000100",
                                4715 => "0000010000",
                                4716 => "0000001000",
                                4717 => "1001110000",
                                4718 => "1011011000",
                                4719 => "1101000000",
                                4720 => "0001011100",
                                4721 => "0100101100",
                                4722 => "0000100100",
                                4723 => "0110000000",
                                4724 => "0011001000",
                                4725 => "1011000100",
                                4726 => "1000110000",
                                4727 => "0100011100",
                                4728 => "0100111100",
                                4729 => "0000100000",
                                4730 => "0000000000",
                                4731 => "0100010101",
                                4732 => "0100010110",
                                4733 => "0000000000",
                                4734 => "0000000000",
                                4735 => "0011000000",
                                4736 => "0000000000",
                                4737 => "0000000000",
                                4738 => "0100000000",
                                4739 => "0000000000",
                                4740 => "1110101100",
                                4741 => "0000011000",
                                4742 => "1110011100",
                                4743 => "1001101100",
                                4744 => "0011011000",
                                4745 => "0101000100",
                                4746 => "1010111100",
                                4747 => "1100110000",
                                4748 => "1100000000",
                                4749 => "1010100000",
                                4750 => "0000000100",
                                4751 => "0110011000",
                                4752 => "0000000100",
                                4753 => "1011101100",
                                4754 => "1110010100",
                                4755 => "0000110100",
                                4756 => "1010111100",
                                4757 => "1000001000",
                                4758 => "1001111000",
                                4759 => "0110001100",
                                4760 => "1010111000",
                                4761 => "1011110000",
                                4762 => "1011000100",
                                4763 => "0000001100",
                                4764 => "0111000000",
                                4765 => "0001001000",
                                4766 => "0110100100",
                                4767 => "0000001100",
                                4768 => "1101110100",
                                4769 => "0111000000",
                                4770 => "0000000000",
                                4771 => "0000000000",
                                4772 => "0000001000",
                                4773 => "0000010000",
                                4774 => "0000010100",
                                4775 => "1011010000",
                                4776 => "0000000100",
                                4777 => "0000000100",
                                4778 => "0000010000",
                                4779 => "0000001000",
                                4780 => "1001110000",
                                4781 => "1011011000",
                                4782 => "1101000000",
                                4783 => "0001011100",
                                4784 => "0100101100",
                                4785 => "0000100100",
                                4786 => "0110000000",
                                4787 => "0011001000",
                                4788 => "1011000100",
                                4789 => "1000110000",
                                4790 => "0100011100",
                                4791 => "0100111100",
                                4792 => "0000100000",
                                4793 => "0000000000",
                                4794 => "0100010101",
                                4795 => "0100010110",
                                4796 => "0000000000",
                                4797 => "0000000000",
                                4798 => "0011000000",
                                4799 => "0000000000",
                                4800 => "0000000000",
                                4801 => "0100000000",
                                4802 => "0000000000",
                                4803 => "1110010000",
                                4804 => "0000011000",
                                4805 => "0111001100",
                                4806 => "1100010100",
                                4807 => "0011111100",
                                4808 => "0010000000",
                                4809 => "0010000100",
                                4810 => "1101010000",
                                4811 => "1100000000",
                                4812 => "1010100000",
                                4813 => "0000000100",
                                4814 => "0110011000",
                                4815 => "0000000100",
                                4816 => "1011101100",
                                4817 => "1110010100",
                                4818 => "0000111000",
                                4819 => "0111101100",
                                4820 => "1100011000",
                                4821 => "1111011100",
                                4822 => "0111000000",
                                4823 => "0111100100",
                                4824 => "1001100000",
                                4825 => "0100000000",
                                4826 => "0111001100",
                                4827 => "0111000000",
                                4828 => "0001001000",
                                4829 => "0110100100",
                                4830 => "0000001100",
                                4831 => "1110001000",
                                4832 => "1111110000",
                                4833 => "0000000000",
                                4834 => "0000000000",
                                4835 => "0000001000",
                                4836 => "0000010000",
                                4837 => "0000010100",
                                4838 => "1011010000",
                                4839 => "0000000100",
                                4840 => "0000000100",
                                4841 => "0000010000",
                                4842 => "0000001000",
                                4843 => "1001110000",
                                4844 => "1011011000",
                                4845 => "1101000000",
                                4846 => "0001011100",
                                4847 => "0100101100",
                                4848 => "0000100100",
                                4849 => "0110000000",
                                4850 => "0011001000",
                                4851 => "1011000100",
                                4852 => "1000110000",
                                4853 => "0100011100",
                                4854 => "0100111100",
                                4855 => "0000100000",
                                4856 => "0000000000",
                                4857 => "0100010101",
                                4858 => "0100010110",
                                4859 => "0000000000",
                                4860 => "0000000000",
                                4861 => "0011000000",
                                4862 => "0000000000",
                                4863 => "0000000000",
                                4864 => "0100000000",
                                4865 => "0000000000",
                                4866 => "1110010100",
                                4867 => "0000011000",
                                4868 => "0111001000",
                                4869 => "1100010100",
                                4870 => "0011111100",
                                4871 => "0010000000",
                                4872 => "0010000100",
                                4873 => "1101010000",
                                4874 => "1100000000",
                                4875 => "1010100000",
                                4876 => "0000000100",
                                4877 => "0110011000",
                                4878 => "0000000100",
                                4879 => "1011101100",
                                4880 => "1110010100",
                                4881 => "0000111100",
                                4882 => "1011100100",
                                4883 => "1101110000",
                                4884 => "0111010100",
                                4885 => "0100001000",
                                4886 => "1110000100",
                                4887 => "0100110100",
                                4888 => "1010011000",
                                4889 => "1001111000",
                                4890 => "0111000000",
                                4891 => "0001001000",
                                4892 => "0110100100",
                                4893 => "0000001100",
                                4894 => "0101100100",
                                4895 => "0011001100",
                                4896 => "0000000000",
                                4897 => "0000000000",
                                4898 => "0000001000",
                                4899 => "0000010000",
                                4900 => "0000010100",
                                4901 => "1011010000",
                                4902 => "0000000100",
                                4903 => "0000000100",
                                4904 => "0000010000",
                                4905 => "0000001000",
                                4906 => "1001110000",
                                4907 => "1011011000",
                                4908 => "1101000000",
                                4909 => "0001011100",
                                4910 => "0100101100",
                                4911 => "0000100100",
                                4912 => "0110000000",
                                4913 => "0011001000",
                                4914 => "1011000100",
                                4915 => "1000110000",
                                4916 => "0100011100",
                                4917 => "0100111100",
                                4918 => "0000100000",
                                4919 => "0000000000",
                                4920 => "0100010101",
                                4921 => "0100010110",
                                4922 => "0000000000",
                                4923 => "0000000000",
                                4924 => "0011000000",
                                4925 => "0001010100",
                                4926 => "0000011000",
                                4927 => "0000000000",
                                4928 => "0000000000",
                                4929 => "1111010000",
                                4930 => "0000011000",
                                4931 => "0100101000",
                                4932 => "0001110100",
                                4933 => "0000110100",
                                4934 => "0010000100",
                                4935 => "1001100000",
                                4936 => "0111010100",
                                4937 => "1100000000",
                                4938 => "1010100000",
                                4939 => "0000000100",
                                4940 => "0110011000",
                                4941 => "0000000100",
                                4942 => "1011101100",
                                4943 => "1110010100",
                                4944 => "0001000000",
                                4945 => "1010000000",
                                4946 => "0111110100",
                                4947 => "1100000100",
                                4948 => "0101010100",
                                4949 => "1110001100",
                                4950 => "1111111000",
                                4951 => "1101101100",
                                4952 => "0010000100",
                                4953 => "0111000000",
                                4954 => "0001001000",
                                4955 => "0000010100",
                                4956 => "1010000000",
                                4957 => "0000111000",
                                4958 => "0001111100",
                                4959 => "0000000000",
                                4960 => "0000000000",
                                4961 => "0000001000",
                                4962 => "0000010000",
                                4963 => "0000010100",
                                4964 => "1010000000",
                                4965 => "0000000100",
                                4966 => "0000000100",
                                4967 => "0000010000",
                                4968 => "0000001000",
                                4969 => "1001110000",
                                4970 => "1011011000",
                                4971 => "1101000000",
                                4972 => "0001011100",
                                4973 => "0100101100",
                                4974 => "0000100100",
                                4975 => "0110000000",
                                4976 => "0011001000",
                                4977 => "1011000100",
                                4978 => "1000110000",
                                4979 => "0100011100",
                                4980 => "0100111100",
                                4981 => "0000100000",
                                4982 => "0000000000",
                                4983 => "0100010101",
                                4984 => "0100010110",
                                4985 => "0000000000",
                                4986 => "0000000000",
                                4987 => "0011000000",
                                4988 => "0001010100",
                                4989 => "0000100000",
                                4990 => "0000000000",
                                4991 => "0000000000",
                                4992 => "1111010000",
                                4993 => "0000011000",
                                4994 => "0100101000",
                                4995 => "0001101100",
                                4996 => "0000110100",
                                4997 => "0010000100",
                                4998 => "1001100000",
                                4999 => "0111010100",
                                5000 => "1100000000",
                                5001 => "1010100000",
                                5002 => "0000000100",
                                5003 => "0110011000",
                                5004 => "0000000100",
                                5005 => "1011101100",
                                5006 => "1110010100",
                                5007 => "0001000000",
                                5008 => "1010000000",
                                5009 => "0111110100",
                                5010 => "1100000100",
                                5011 => "0101010100",
                                5012 => "1110001100",
                                5013 => "1111111000",
                                5014 => "1101101100",
                                5015 => "0010000100",
                                5016 => "0111000000",
                                5017 => "0001001000",
                                5018 => "0000010100",
                                5019 => "1010000000",
                                5020 => "0000111000",
                                5021 => "0001111100",
                                5022 => "0000000000",
                                5023 => "0000000000",
                                5024 => "0000001000",
                                5025 => "0000010000",
                                5026 => "0000010100",
                                5027 => "1010000000",
                                5028 => "0000000100",
                                5029 => "0000000100",
                                5030 => "0000010000",
                                5031 => "0000001000",
                                5032 => "1001110000",
                                5033 => "1011011000",
                                5034 => "1101000000",
                                5035 => "0001011100",
                                5036 => "0100101100",
                                5037 => "0000100100",
                                5038 => "0110000000",
                                5039 => "0011001000",
                                5040 => "1011000100",
                                5041 => "1000110000",
                                5042 => "0100011100",
                                5043 => "0100111100",
                                5044 => "0000100000",
                                5045 => "0000000000",
                                5046 => "0100010101",
                                5047 => "0100010110",
                                5048 => "0000000000",
                                5049 => "0000000000",
                                5050 => "0011000000",
                                5051 => "0100101000",
                                5052 => "1000101000",
                                5053 => "0100000000",
                                5054 => "0000000000",
                                5055 => "1111000000",
                                5056 => "0000011000",
                                5057 => "0110100100",
                                5058 => "1110001100",
                                5059 => "1100000000",
                                5060 => "0010011000",
                                5061 => "0101010000",
                                5062 => "0010010100",
                                5063 => "1100000000",
                                5064 => "1010100000",
                                5065 => "0000000100",
                                5066 => "0110011000",
                                5067 => "0000000100",
                                5068 => "1011101100",
                                5069 => "1110010100",
                                5070 => "0001000100",
                                5071 => "1111000100",
                                5072 => "0100100000",
                                5073 => "1111101100",
                                5074 => "1100110000",
                                5075 => "0101001100",
                                5076 => "0110111100",
                                5077 => "0011110000",
                                5078 => "1010010100",
                                5079 => "0111000000",
                                5080 => "0001001000",
                                5081 => "0011100100",
                                5082 => "0000100000",
                                5083 => "0001000000",
                                5084 => "1011011100",
                                5085 => "0000000000",
                                5086 => "0000000000",
                                5087 => "0000001000",
                                5088 => "0000010000",
                                5089 => "0000010100",
                                5090 => "1011010000",
                                5091 => "0000010000",
                                5092 => "0000001000",
                                5093 => "0000000000",
                                5094 => "0000000000",
                                5095 => "1001110000",
                                5096 => "1011011000",
                                5097 => "1101000000",
                                5098 => "0001011100",
                                5099 => "0100101100",
                                5100 => "0000100100",
                                5101 => "0110000000",
                                5102 => "0011001000",
                                5103 => "1011000100",
                                5104 => "1000110000",
                                5105 => "0100011100",
                                5106 => "0100111100",
                                5107 => "0000100000",
                                5108 => "0000000000",
                                5109 => "0100010101",
                                5110 => "0100010110",
                                5111 => "0000000000",
                                5112 => "0000000000",
                                5113 => "0011000000",
                                5114 => "0000000000",
                                5115 => "0000000000",
                                5116 => "0100000000",
                                5117 => "0000000000",
                                5118 => "0011000100",
                                5119 => "0000011000",
                                5120 => "1000100100",
                                5121 => "0100110100",
                                5122 => "1000110000",
                                5123 => "0101001000",
                                5124 => "0111001000",
                                5125 => "0001101000",
                                5126 => "1100000000",
                                5127 => "1010100000",
                                5128 => "0000000100",
                                5129 => "0110011000",
                                5130 => "0000000100",
                                5131 => "1011101100",
                                5132 => "1110010100",
                                5133 => "0001001000",
                                5134 => "0001010000",
                                5135 => "1011001100",
                                5136 => "1001100000",
                                5137 => "1010100000",
                                5138 => "1111010100",
                                5139 => "0100001000",
                                5140 => "1011111100",
                                5141 => "1001001000",
                                5142 => "0111000000",
                                5143 => "0001001000",
                                5144 => "1111111100",
                                5145 => "1111111100",
                                5146 => "0111100100",
                                5147 => "1010110100",
                                5148 => "0000000000",
                                5149 => "0000000000",
                                5150 => "0000001000",
                                5151 => "0000010000",
                                5152 => "0000010100",
                                5153 => "1001110000",
                                5154 => "0000000100",
                                5155 => "0000000100",
                                5156 => "0000010000",
                                5157 => "0000001000",
                                5158 => "1001110000",
                                5159 => "1011011000",
                                5160 => "1101000000",
                                5161 => "0001011100",
                                5162 => "0100101100",
                                5163 => "0000100100",
                                5164 => "0110000000",
                                5165 => "0011001000",
                                5166 => "1011000100",
                                5167 => "1000110000",
                                5168 => "0100011100",
                                5169 => "0100111100",
                                5170 => "0000100000",
                                5171 => "0000000000",
                                5172 => "0100010101",
                                5173 => "0100010110",
                                5174 => "0000000000",
                                5175 => "0000000000",
                                5176 => "0011000000",
                                5177 => "0111001000",
                                5178 => "0111000000",
                                5179 => "0100000000",
                                5180 => "0000000000",
                                5181 => "1110111100",
                                5182 => "0000011000",
                                5183 => "0100001000",
                                5184 => "1111110100",
                                5185 => "1100000000",
                                5186 => "0010011000",
                                5187 => "0101010000",
                                5188 => "0010010100",
                                5189 => "1100000000",
                                5190 => "1010100000",
                                5191 => "0000000100",
                                5192 => "0110011000",
                                5193 => "0000000100",
                                5194 => "1011101100",
                                5195 => "1110010100",
                                5196 => "0001001100",
                                5197 => "1101011100",
                                5198 => "1011001000",
                                5199 => "1001010000",
                                5200 => "0110110000",
                                5201 => "0111010000",
                                5202 => "0110011100",
                                5203 => "0100101100",
                                5204 => "0100001000",
                                5205 => "0111000000",
                                5206 => "0001001000",
                                5207 => "0011100100",
                                5208 => "0000100000",
                                5209 => "0110001000",
                                5210 => "0001011000",
                                5211 => "0000000000",
                                5212 => "0000000000",
                                5213 => "0000001000",
                                5214 => "0000010000",
                                5215 => "0000010100",
                                5216 => "1011010000",
                                5217 => "0000010000",
                                5218 => "0000001000",
                                5219 => "0000000000",
                                5220 => "0000000000",
                                5221 => "1001110000",
                                5222 => "1011011000",
                                5223 => "1101000000",
                                5224 => "0001011100",
                                5225 => "0100101100",
                                5226 => "0000100100",
                                5227 => "0110000000",
                                5228 => "0011001000",
                                5229 => "1011000100",
                                5230 => "1000110000",
                                5231 => "0100011100",
                                5232 => "0100111100",
                                5233 => "0000100000",
                                5234 => "0000000000",
                                5235 => "0100010101",
                                5236 => "0100010110",
                                5237 => "0000000000",
                                5238 => "0000000000",
                                5239 => "0011000000",
                                5240 => "0000000000",
                                5241 => "0000000000",
                                5242 => "0100000000",
                                5243 => "0000000000",
                                5244 => "0011100000",
                                5245 => "0000011000",
                                5246 => "1000110100",
                                5247 => "1111100000",
                                5248 => "1100011100",
                                5249 => "1110100000",
                                5250 => "0010101000",
                                5251 => "1101100100",
                                5252 => "1100000000",
                                5253 => "1010100000",
                                5254 => "0000000100",
                                5255 => "0110011000",
                                5256 => "0000000100",
                                5257 => "1011101100",
                                5258 => "1110010100",
                                5259 => "0001010000",
                                5260 => "0110101100",
                                5261 => "0001011100",
                                5262 => "0000101000",
                                5263 => "0011000100",
                                5264 => "1100100100",
                                5265 => "0110101100",
                                5266 => "1000101100",
                                5267 => "1101110100",
                                5268 => "0111000000",
                                5269 => "0001001000",
                                5270 => "1111111100",
                                5271 => "1111111100",
                                5272 => "0001110000",
                                5273 => "1101111000",
                                5274 => "0000000000",
                                5275 => "0000000000",
                                5276 => "0000001000",
                                5277 => "0000010000",
                                5278 => "0000010100",
                                5279 => "1011010000",
                                5280 => "0000000100",
                                5281 => "0000000100",
                                5282 => "0000010000",
                                5283 => "0000001000",
                                5284 => "1001110000",
                                5285 => "1011011000",
                                5286 => "1101000000",
                                5287 => "0001011100",
                                5288 => "0100101100",
                                5289 => "0000100100",
                                5290 => "0110000000",
                                5291 => "0011001000",
                                5292 => "1011000100",
                                5293 => "1000110000",
                                5294 => "0100011100",
                                5295 => "0100111100",
                                5296 => "0000100000",
                                5297 => "0000000000",
                                5298 => "0100010101",
                                5299 => "0100010110",
                                5300 => "0000000000",
                                5301 => "0000000000",
                                5302 => "0011000000",
                                5303 => "0000000000",
                                5304 => "0000000000",
                                5305 => "0100000000",
                                5306 => "0000000000",
                                5307 => "0011001100",
                                5308 => "0000011000",
                                5309 => "1000000000",
                                5310 => "0110001000",
                                5311 => "1000110000",
                                5312 => "0101001000",
                                5313 => "0111100100",
                                5314 => "0000010100",
                                5315 => "1100000000",
                                5316 => "1010100000",
                                5317 => "0000000100",
                                5318 => "0110011000",
                                5319 => "0000000100",
                                5320 => "1011101100",
                                5321 => "1110010100",
                                5322 => "0001010100",
                                5323 => "1111100100",
                                5324 => "1001110000",
                                5325 => "1000011100",
                                5326 => "1110100100",
                                5327 => "0000110000",
                                5328 => "0100110000",
                                5329 => "0000011000",
                                5330 => "0000010000",
                                5331 => "0111000000",
                                5332 => "0001001000",
                                5333 => "1111111100",
                                5334 => "1111111100",
                                5335 => "0100000100",
                                5336 => "0001101000",
                                5337 => "0000000000",
                                5338 => "0000000000",
                                5339 => "0000001000",
                                5340 => "0000010000",
                                5341 => "0000010100",
                                5342 => "1001110000",
                                5343 => "0000000100",
                                5344 => "0000000100",
                                5345 => "0000010000",
                                5346 => "0000001000",
                                5347 => "1001110000",
                                5348 => "1011011000",
                                5349 => "1101000000",
                                5350 => "0001011100",
                                5351 => "0100101100",
                                5352 => "0000100100",
                                5353 => "0110000000",
                                5354 => "0011001000",
                                5355 => "1011000100",
                                5356 => "1000110000",
                                5357 => "0100011100",
                                5358 => "0100111100",
                                5359 => "0000100000",
                                5360 => "0000000000",
                                5361 => "0100010101",
                                5362 => "0100010110",
                                5363 => "0000000000",
                                5364 => "0000000000",
                                5365 => "0011000000",
                                5366 => "1010011000",
                                5367 => "1011000000",
                                5368 => "0100000000",
                                5369 => "0000000000",
                                5370 => "1110111100",
                                5371 => "0000011000",
                                5372 => "0000111000",
                                5373 => "1011110100",
                                5374 => "1100000000",
                                5375 => "0010011000",
                                5376 => "0101010000",
                                5377 => "0010010100",
                                5378 => "1100000000",
                                5379 => "1010100000",
                                5380 => "0000000100",
                                5381 => "0110011000",
                                5382 => "0000000100",
                                5383 => "1011101100",
                                5384 => "1110010100",
                                5385 => "0001011000",
                                5386 => "1101000000",
                                5387 => "1001111100",
                                5388 => "0010001100",
                                5389 => "0011110100",
                                5390 => "0111001100",
                                5391 => "1101011100",
                                5392 => "1100111000",
                                5393 => "0001101100",
                                5394 => "0111000000",
                                5395 => "0001001000",
                                5396 => "0011100100",
                                5397 => "0000100000",
                                5398 => "0101100000",
                                5399 => "0000110000",
                                5400 => "0000000000",
                                5401 => "0000000000",
                                5402 => "0000001000",
                                5403 => "0000010000",
                                5404 => "0000010100",
                                5405 => "1011010000",
                                5406 => "0000010000",
                                5407 => "0000001000",
                                5408 => "0000000000",
                                5409 => "0000000000",
                                5410 => "1001110000",
                                5411 => "1011011000",
                                5412 => "1101000000",
                                5413 => "0001011100",
                                5414 => "0100101100",
                                5415 => "0000100100",
                                5416 => "0110000000",
                                5417 => "0011001000",
                                5418 => "1011000100",
                                5419 => "1000110000",
                                5420 => "0100011100",
                                5421 => "0100111100",
                                5422 => "0000100000",
                                5423 => "0000000000",
                                5424 => "0100010101",
                                5425 => "0100010110",
                                5426 => "0000000000",
                                5427 => "0000000000",
                                5428 => "0011000000",
                                5429 => "0000000000",
                                5430 => "0000000000",
                                5431 => "0100000000",
                                5432 => "0000000000",
                                5433 => "0011010100",
                                5434 => "0000011000",
                                5435 => "0001011000",
                                5436 => "1101010000",
                                5437 => "0110100000",
                                5438 => "0001101000",
                                5439 => "0000010000",
                                5440 => "1100110000",
                                5441 => "1100000000",
                                5442 => "1010100000",
                                5443 => "0000000100",
                                5444 => "0110011000",
                                5445 => "0000000100",
                                5446 => "1011101100",
                                5447 => "1110010100",
                                5448 => "0001011100",
                                5449 => "0101011000",
                                5450 => "1111000000",
                                5451 => "1100101100",
                                5452 => "1010101000",
                                5453 => "0001011000",
                                5454 => "1000001100",
                                5455 => "1000101000",
                                5456 => "0001111000",
                                5457 => "0111000000",
                                5458 => "0001001000",
                                5459 => "1111111100",
                                5460 => "1111111100",
                                5461 => "1010101000",
                                5462 => "0100011100",
                                5463 => "0000000000",
                                5464 => "0000000000",
                                5465 => "0000001000",
                                5466 => "0000010000",
                                5467 => "0000010100",
                                5468 => "0111100000",
                                5469 => "0000000100",
                                5470 => "0000000100",
                                5471 => "0000010000",
                                5472 => "0000001000",
                                5473 => "1001110000",
                                5474 => "1011011000",
                                5475 => "1101000000",
                                5476 => "0001011100",
                                5477 => "0100101100",
                                5478 => "0000100100",
                                5479 => "0110000000",
                                5480 => "0011001000",
                                5481 => "1011000100",
                                5482 => "1000110000",
                                5483 => "0100011100",
                                5484 => "0100111100",
                                5485 => "0000100000",
                                5486 => "0000000000",
                                5487 => "0100010101",
                                5488 => "0100010110",
                                5489 => "0000000000",
                                5490 => "0000000000",
                                5491 => "0011000000",
                                5492 => "0101011000",
                                5493 => "1001101100",
                                5494 => "0000000000",
                                5495 => "0000000000",
                                5496 => "1111010000",
                                5497 => "0000011000",
                                5498 => "0000100000",
                                5499 => "1000100000",
                                5500 => "0000110100",
                                5501 => "0010000100",
                                5502 => "1001100000",
                                5503 => "0111010100",
                                5504 => "1100000000",
                                5505 => "1010100000",
                                5506 => "0000000100",
                                5507 => "0110011000",
                                5508 => "0000000100",
                                5509 => "1011101100",
                                5510 => "1110010100",
                                5511 => "0001100000",
                                5512 => "1111111100",
                                5513 => "0011100000",
                                5514 => "1010100100",
                                5515 => "0110001100",
                                5516 => "1110010000",
                                5517 => "0101001100",
                                5518 => "1000010000",
                                5519 => "0111000100",
                                5520 => "0111000000",
                                5521 => "0001001000",
                                5522 => "0000010100",
                                5523 => "1010000000",
                                5524 => "0001110100",
                                5525 => "1010100100",
                                5526 => "0000000000",
                                5527 => "0000000000",
                                5528 => "0000001000",
                                5529 => "0000010000",
                                5530 => "0000010100",
                                5531 => "1010000000",
                                5532 => "0000000100",
                                5533 => "0000000100",
                                5534 => "0000010000",
                                5535 => "0000001000",
                                5536 => "1001110000",
                                5537 => "1011011000",
                                5538 => "1101000000",
                                5539 => "0001011100",
                                5540 => "0100101100",
                                5541 => "0000100100",
                                5542 => "0110000000",
                                5543 => "0011001000",
                                5544 => "1011000100",
                                5545 => "1000110000",
                                5546 => "0100011100",
                                5547 => "0100111100",
                                5548 => "0000100000",
                                5549 => "0000000000",
                                5550 => "0100010101",
                                5551 => "0100010110",
                                5552 => "0000000000",
                                5553 => "0000000000",
                                5554 => "0011000000",
                                5555 => "0000010100",
                                5556 => "1010100000",
                                5557 => "0000000000",
                                5558 => "0000000000",
                                5559 => "1111001100",
                                5560 => "0000011000",
                                5561 => "0110011100",
                                5562 => "1110001100",
                                5563 => "0000110100",
                                5564 => "0010000100",
                                5565 => "1000101100",
                                5566 => "0000110100",
                                5567 => "1100000000",
                                5568 => "1010100000",
                                5569 => "0000000100",
                                5570 => "0110011000",
                                5571 => "0000000100",
                                5572 => "1011101100",
                                5573 => "1110010100",
                                5574 => "0001100100",
                                5575 => "1100101000",
                                5576 => "0011011100",
                                5577 => "1010010000",
                                5578 => "0101100100",
                                5579 => "1011010100",
                                5580 => "0101001100",
                                5581 => "0110100100",
                                5582 => "0011101000",
                                5583 => "0111000000",
                                5584 => "0001001000",
                                5585 => "0000010100",
                                5586 => "1010000000",
                                5587 => "1010111100",
                                5588 => "0101001000",
                                5589 => "0000000000",
                                5590 => "0000000000",
                                5591 => "0000001000",
                                5592 => "0000010000",
                                5593 => "0000010100",
                                5594 => "1010000000",
                                5595 => "0000000100",
                                5596 => "0000000100",
                                5597 => "0000010000",
                                5598 => "0000001000",
                                5599 => "0000001000");
    
    
   begin
    data_out <= ROM(to_integer(unsigned(unsigned(address))));
  end architecture;
