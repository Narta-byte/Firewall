--Hello i am a file