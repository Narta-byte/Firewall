-- cecil
