--this is a test file