LIBRARY IEEE;
LIBRARY std;
USE IEEE.std_logic_1164.ALL;
--USE IEEE.numeric_std_unsigned.ALL;
--USE IEEE.numeric_std_unsigned;
USE IEEE.NUMERIC_STD.ALL;

ENTITY INPUT_ROM IS
PORT (
    address : IN STD_LOGIC_VECTOR(15 DOWNTO 0); --64 addresses
    data_out : OUT STD_LOGIC_VECTOR(8 DOWNTO 0) --9 bits, the lsb is start_of_data, and the 8 others are the ip header
);
END ENTITY;

ARCHITECTURE INPUT_ROM_arch OF INPUT_ROM IS
 type ROM_type is array (0 to 9707) of std_logic_vector(8 downto 0);

constant ROM : ROM_type := (0 => "000000000",
                            1 => "000000000",
                            2 => "000011000",
                            3 => "100111110",
                            4 => "111100100",
                            5 => "010101110",
                            6 => "100111000",
                            7 => "101101100",
                            8 => "110100000",
                            9 => "000101110",
                            10 => "010010110",
                            11 => "000010010",
                            12 => "000010000",
                            13 => "000000000",
                            14 => "010001011",
                            15 => "100110000",
                            16 => "000000000",
                            17 => "010001010",
                            18 => "111100100",
                            19 => "011001100",
                            20 => "010000000",
                            21 => "000000000",
                            22 => "100000000",
                            23 => "000001100",
                            24 => "101000000",
                            25 => "010101000",
                            26 => "000010100",
                            27 => "110100010",
                            28 => "111101010",
                            29 => "011010110",
                            30 => "000111110",
                            31 => "000011010",
                            32 => "010010000",
                            33 => "000101100",
                            34 => "111001110",
                            35 => "001010100",
                            36 => "000000010",
                            37 => "101110110",
                            38 => "000011100",
                            39 => "101000100",
                            40 => "011110000",
                            41 => "110010100",
                            42 => "110100000",
                            43 => "001010110",
                            44 => "001010010",
                            45 => "100110010",
                            46 => "010100000",
                            47 => "000110000",
                            48 => "000000010",
                            49 => "111111110",
                            50 => "011110100",
                            51 => "110111010",
                            52 => "000000000",
                            53 => "000000000",
                            54 => "000101110",
                            55 => "000000110",
                            56 => "000000110",
                            57 => "000000000",
                            58 => "000110000",
                            59 => "111100010",
                            60 => "001110100",
                            61 => "110000010",
                            62 => "111100010",
                            63 => "110010000",
                            64 => "110110000",
                            65 => "110010010",
                            66 => "010001000",
                            67 => "110001010",
                            68 => "100001010",
                            69 => "001100010",
                            70 => "001011100",
                            71 => "110110000",
                            72 => "110011100",
                            73 => "111111100",
                            74 => "011010110",
                            75 => "010010010",
                            76 => "001000000",
                            77 => "000100010",
                            78 => "101100110",
                            79 => "101001110",
                            80 => "110010010",
                            81 => "010000110",
                            82 => "010110010",
                            83 => "000000000",
                            84 => "000000000",
                            85 => "000011000",
                            86 => "100111110",
                            87 => "111100100",
                            88 => "010101110",
                            89 => "100111000",
                            90 => "101101100",
                            91 => "110100000",
                            92 => "000101110",
                            93 => "010010110",
                            94 => "000010010",
                            95 => "000010000",
                            96 => "000000000",
                            97 => "010001011",
                            98 => "100110000",
                            99 => "000000000",
                            100 => "010001010",
                            101 => "111100100",
                            102 => "011001110",
                            103 => "010000000",
                            104 => "000000000",
                            105 => "100000000",
                            106 => "000001100",
                            107 => "101000000",
                            108 => "010100110",
                            109 => "000010100",
                            110 => "110100010",
                            111 => "111101010",
                            112 => "011010110",
                            113 => "000111110",
                            114 => "000011010",
                            115 => "010010000",
                            116 => "000101100",
                            117 => "110011000",
                            118 => "000110110",
                            119 => "000000010",
                            120 => "101110110",
                            121 => "011111110",
                            122 => "011100100",
                            123 => "011011010",
                            124 => "100010110",
                            125 => "111110000",
                            126 => "101011010",
                            127 => "111011000",
                            128 => "011101010",
                            129 => "010100000",
                            130 => "000110000",
                            131 => "000000010",
                            132 => "111111010",
                            133 => "100000010",
                            134 => "000001010",
                            135 => "000000000",
                            136 => "000000000",
                            137 => "000101110",
                            138 => "000000110",
                            139 => "000000110",
                            140 => "000000000",
                            141 => "000110000",
                            142 => "100010010",
                            143 => "001000110",
                            144 => "110101010",
                            145 => "101100000",
                            146 => "011110100",
                            147 => "110101000",
                            148 => "000111110",
                            149 => "111101110",
                            150 => "011010000",
                            151 => "001111000",
                            152 => "010111010",
                            153 => "000101000",
                            154 => "000000010",
                            155 => "101010100",
                            156 => "000010100",
                            157 => "100110100",
                            158 => "000000000",
                            159 => "000000110",
                            160 => "101000000",
                            161 => "000000100",
                            162 => "011011100",
                            163 => "010000110",
                            164 => "011110000",
                            165 => "011101010",
                            166 => "000000000",
                            167 => "000000000",
                            168 => "000011000",
                            169 => "100111110",
                            170 => "111100100",
                            171 => "010101110",
                            172 => "100111000",
                            173 => "101101100",
                            174 => "110100000",
                            175 => "000101110",
                            176 => "010010110",
                            177 => "000010010",
                            178 => "000010000",
                            179 => "000000000",
                            180 => "010001011",
                            181 => "100110000",
                            182 => "000000000",
                            183 => "010001010",
                            184 => "111100100",
                            185 => "011010000",
                            186 => "010000000",
                            187 => "000000000",
                            188 => "100000000",
                            189 => "000001100",
                            190 => "101000000",
                            191 => "010100100",
                            192 => "000010100",
                            193 => "110100010",
                            194 => "111101010",
                            195 => "011010110",
                            196 => "000111110",
                            197 => "000011010",
                            198 => "010010000",
                            199 => "000101100",
                            200 => "111001110",
                            201 => "001011000",
                            202 => "000000010",
                            203 => "101110110",
                            204 => "101000110",
                            205 => "011100100",
                            206 => "001000100",
                            207 => "000100100",
                            208 => "111110010",
                            209 => "001110000",
                            210 => "010000100",
                            211 => "100000100",
                            212 => "010100000",
                            213 => "000110000",
                            214 => "000000100",
                            215 => "000000000",
                            216 => "100011100",
                            217 => "000110100",
                            218 => "000000000",
                            219 => "000000000",
                            220 => "000101110",
                            221 => "000000110",
                            222 => "000000110",
                            223 => "000000000",
                            224 => "000110000",
                            225 => "001000110",
                            226 => "101100010",
                            227 => "110100000",
                            228 => "011111000",
                            229 => "011101100",
                            230 => "000010110",
                            231 => "010011100",
                            232 => "000000000",
                            233 => "010100100",
                            234 => "011100100",
                            235 => "010111100",
                            236 => "111001010",
                            237 => "100110110",
                            238 => "000111110",
                            239 => "100101110",
                            240 => "111110000",
                            241 => "111111010",
                            242 => "011011110",
                            243 => "010101110",
                            244 => "110110010",
                            245 => "100111100",
                            246 => "001001010",
                            247 => "011110100",
                            248 => "100000110",
                            249 => "000000000",
                            250 => "000000000",
                            251 => "000011000",
                            252 => "100111110",
                            253 => "111100100",
                            254 => "010101110",
                            255 => "100111000",
                            256 => "101101100",
                            257 => "110100000",
                            258 => "000101110",
                            259 => "010010110",
                            260 => "000010010",
                            261 => "000010000",
                            262 => "000000000",
                            263 => "010001011",
                            264 => "100110000",
                            265 => "000000000",
                            266 => "010001010",
                            267 => "111100100",
                            268 => "011010010",
                            269 => "010000000",
                            270 => "000000000",
                            271 => "100000000",
                            272 => "000001100",
                            273 => "101000000",
                            274 => "010100010",
                            275 => "000010100",
                            276 => "110100010",
                            277 => "111101010",
                            278 => "011010110",
                            279 => "000111110",
                            280 => "000011010",
                            281 => "010010000",
                            282 => "000101100",
                            283 => "111001110",
                            284 => "001010010",
                            285 => "000000010",
                            286 => "101110110",
                            287 => "001100010",
                            288 => "000010100",
                            289 => "110001100",
                            290 => "111000110",
                            291 => "001001010",
                            292 => "111000010",
                            293 => "000111110",
                            294 => "010010010",
                            295 => "010100000",
                            296 => "000110000",
                            297 => "000000100",
                            298 => "000000000",
                            299 => "010000010",
                            300 => "001111110",
                            301 => "000000000",
                            302 => "000000000",
                            303 => "000101110",
                            304 => "000000110",
                            305 => "000000110",
                            306 => "000000000",
                            307 => "000110000",
                            308 => "110010100",
                            309 => "100100000",
                            310 => "011110100",
                            311 => "000111010",
                            312 => "011111000",
                            313 => "111001110",
                            314 => "110010010",
                            315 => "110111010",
                            316 => "101110110",
                            317 => "100110110",
                            318 => "000110010",
                            319 => "011001010",
                            320 => "101001000",
                            321 => "011000010",
                            322 => "101100110",
                            323 => "011011110",
                            324 => "011001010",
                            325 => "100101010",
                            326 => "001101010",
                            327 => "001010110",
                            328 => "101011110",
                            329 => "010111010",
                            330 => "000011100",
                            331 => "010010010",
                            332 => "100111000",
                            333 => "101101100",
                            334 => "110100000",
                            335 => "000101110",
                            336 => "010010110",
                            337 => "000010010",
                            338 => "000000000",
                            339 => "001001110",
                            340 => "100100000",
                            341 => "111001100",
                            342 => "001000010",
                            343 => "010101110",
                            344 => "000010000",
                            345 => "000000000",
                            346 => "010001011",
                            347 => "000000000",
                            348 => "000000000",
                            349 => "011111110",
                            350 => "110111000",
                            351 => "010010100",
                            352 => "010000000",
                            353 => "000000000",
                            354 => "001101000",
                            355 => "000001100",
                            356 => "001111100",
                            357 => "011010000",
                            358 => "101000100",
                            359 => "100111110",
                            360 => "100010000",
                            361 => "111010100",
                            362 => "000010100",
                            363 => "110100010",
                            364 => "111101010",
                            365 => "011010110",
                            366 => "000000010",
                            367 => "101110110",
                            368 => "111001110",
                            369 => "000101110",
                            370 => "000011110",
                            371 => "001010110",
                            372 => "100010010",
                            373 => "101101010",
                            374 => "011101110",
                            375 => "001011010",
                            376 => "101000110",
                            377 => "110001100",
                            378 => "010100000",
                            379 => "000110000",
                            380 => "000000000",
                            381 => "010101000",
                            382 => "100110100",
                            383 => "101010010",
                            384 => "000000000",
                            385 => "000000000",
                            386 => "000101110",
                            387 => "000000110",
                            388 => "000000110",
                            389 => "000000000",
                            390 => "010100100",
                            391 => "001100110",
                            392 => "011010010",
                            393 => "000101110",
                            394 => "001110010",
                            395 => "111110100",
                            396 => "000000000",
                            397 => "001111100",
                            398 => "100100110",
                            399 => "100100100",
                            400 => "100001010",
                            401 => "111100000",
                            402 => "111010010",
                            403 => "001001000",
                            404 => "110111010",
                            405 => "000000100",
                            406 => "000001000",
                            407 => "101100010",
                            408 => "100001100",
                            409 => "101101100",
                            410 => "110010110",
                            411 => "010101110",
                            412 => "000010010",
                            413 => "101100100",
                            414 => "111000000",
                            415 => "011101110",
                            416 => "001110010",
                            417 => "101011000",
                            418 => "011110100",
                            419 => "001011110",
                            420 => "101011010",
                            421 => "100001000",
                            422 => "101001000",
                            423 => "011101110",
                            424 => "110011110",
                            425 => "000010100",
                            426 => "111010000",
                            427 => "000010110",
                            428 => "011101000",
                            429 => "110101000",
                            430 => "011001000",
                            431 => "110111000",
                            432 => "000101010",
                            433 => "111011000",
                            434 => "010010110",
                            435 => "000011010",
                            436 => "101010100",
                            437 => "111110100",
                            438 => "000100010",
                            439 => "000100100",
                            440 => "000111100",
                            441 => "011110100",
                            442 => "011000010",
                            443 => "111000000",
                            444 => "101101000",
                            445 => "101111010",
                            446 => "111111110",
                            447 => "010001010",
                            448 => "001011100",
                            449 => "011011100",
                            450 => "010011110",
                            451 => "001110110",
                            452 => "110111010",
                            453 => "010001000",
                            454 => "000000000",
                            455 => "010010110",
                            456 => "011000100",
                            457 => "110100110",
                            458 => "100000110",
                            459 => "001100000",
                            460 => "111101110",
                            461 => "011000000",
                            462 => "111101000",
                            463 => "100101100",
                            464 => "010011110",
                            465 => "000100000",
                            466 => "111011000",
                            467 => "001001010",
                            468 => "110100110",
                            469 => "100011110",
                            470 => "111101110",
                            471 => "111100000",
                            472 => "000000000",
                            473 => "100111000",
                            474 => "101101100",
                            475 => "110100000",
                            476 => "000101110",
                            477 => "010010110",
                            478 => "000010010",
                            479 => "000000000",
                            480 => "001001110",
                            481 => "100100000",
                            482 => "111001100",
                            483 => "001000010",
                            484 => "010101110",
                            485 => "000010000",
                            486 => "000000000",
                            487 => "010001011",
                            488 => "000000000",
                            489 => "000000000",
                            490 => "001010000",
                            491 => "110100010",
                            492 => "101000110",
                            493 => "010000000",
                            494 => "000000000",
                            495 => "010100100",
                            496 => "000001100",
                            497 => "111011110",
                            498 => "110011000",
                            499 => "000111110",
                            500 => "000011010",
                            501 => "010010000",
                            502 => "000101100",
                            503 => "000010100",
                            504 => "110100010",
                            505 => "111101010",
                            506 => "011010110",
                            507 => "000000010",
                            508 => "101110110",
                            509 => "111001110",
                            510 => "001010100",
                            511 => "110100000",
                            512 => "001010110",
                            513 => "001010010",
                            514 => "100110010",
                            515 => "000011100",
                            516 => "101000100",
                            517 => "011110000",
                            518 => "111001110",
                            519 => "010100000",
                            520 => "000100000",
                            521 => "000001000",
                            522 => "010010100",
                            523 => "110110010",
                            524 => "111101100",
                            525 => "000000000",
                            526 => "000000000",
                            527 => "100111000",
                            528 => "101101100",
                            529 => "110100000",
                            530 => "000101110",
                            531 => "010010110",
                            532 => "000010010",
                            533 => "000000000",
                            534 => "001001110",
                            535 => "100100000",
                            536 => "111001100",
                            537 => "001000010",
                            538 => "010101110",
                            539 => "000010000",
                            540 => "000000000",
                            541 => "010001011",
                            542 => "000000000",
                            543 => "000000000",
                            544 => "001010000",
                            545 => "101001100",
                            546 => "101111100",
                            547 => "010000000",
                            548 => "000000000",
                            549 => "010100010",
                            550 => "000001100",
                            551 => "000110110",
                            552 => "101100100",
                            553 => "000111110",
                            554 => "000011010",
                            555 => "010010000",
                            556 => "000101100",
                            557 => "000010100",
                            558 => "110100010",
                            559 => "111101010",
                            560 => "011010110",
                            561 => "000000010",
                            562 => "101110110",
                            563 => "110011000",
                            564 => "000110110",
                            565 => "111110000",
                            566 => "101011010",
                            567 => "111011000",
                            568 => "011101010",
                            569 => "011111110",
                            570 => "011100100",
                            571 => "011011010",
                            572 => "101010000",
                            573 => "010100000",
                            574 => "000100000",
                            575 => "000000010",
                            576 => "101001100",
                            577 => "101001100",
                            578 => "101110010",
                            579 => "000000000",
                            580 => "000000000",
                            581 => "100111000",
                            582 => "101101100",
                            583 => "110100000",
                            584 => "000101110",
                            585 => "010010110",
                            586 => "000010010",
                            587 => "000000000",
                            588 => "001001110",
                            589 => "100100000",
                            590 => "111001100",
                            591 => "001000010",
                            592 => "010101110",
                            593 => "000010000",
                            594 => "000000000",
                            595 => "010001011",
                            596 => "000000000",
                            597 => "000000000",
                            598 => "001010000",
                            599 => "001001110",
                            600 => "101110100",
                            601 => "010000000",
                            602 => "000000000",
                            603 => "010100100",
                            604 => "000001100",
                            605 => "100110010",
                            606 => "101101100",
                            607 => "000111110",
                            608 => "000011010",
                            609 => "010010000",
                            610 => "000101100",
                            611 => "000010100",
                            612 => "110100010",
                            613 => "111101010",
                            614 => "011010110",
                            615 => "000000010",
                            616 => "101110110",
                            617 => "111001110",
                            618 => "001010010",
                            619 => "001001010",
                            620 => "111000010",
                            621 => "000111110",
                            622 => "010010010",
                            623 => "001100010",
                            624 => "000010100",
                            625 => "110001110",
                            626 => "000000000",
                            627 => "010100000",
                            628 => "000100000",
                            629 => "000000010",
                            630 => "001001110",
                            631 => "001000010",
                            632 => "001101000",
                            633 => "000000000",
                            634 => "000000000",
                            635 => "100111000",
                            636 => "101101100",
                            637 => "110100000",
                            638 => "000101110",
                            639 => "010010110",
                            640 => "000010010",
                            641 => "000000000",
                            642 => "001001110",
                            643 => "100100000",
                            644 => "111001100",
                            645 => "001000010",
                            646 => "010101110",
                            647 => "000010000",
                            648 => "000000000",
                            649 => "010001011",
                            650 => "000000000",
                            651 => "000000000",
                            652 => "001010000",
                            653 => "010011000",
                            654 => "000110100",
                            655 => "010000000",
                            656 => "000000000",
                            657 => "010100010",
                            658 => "000001100",
                            659 => "011101100",
                            660 => "010101100",
                            661 => "000111110",
                            662 => "000011010",
                            663 => "010010000",
                            664 => "000101100",
                            665 => "000010100",
                            666 => "110100010",
                            667 => "111101010",
                            668 => "011010110",
                            669 => "000000010",
                            670 => "101110110",
                            671 => "111001110",
                            672 => "001011000",
                            673 => "111110010",
                            674 => "001110000",
                            675 => "010000100",
                            676 => "100000100",
                            677 => "101000110",
                            678 => "011100100",
                            679 => "001000100",
                            680 => "001011110",
                            681 => "010100000",
                            682 => "000100000",
                            683 => "000000010",
                            684 => "001011000",
                            685 => "010111010",
                            686 => "000001000",
                            687 => "000000000",
                            688 => "000000000",
                            689 => "100111000",
                            690 => "101101100",
                            691 => "110100000",
                            692 => "000101110",
                            693 => "010010110",
                            694 => "000010010",
                            695 => "000000000",
                            696 => "001001110",
                            697 => "100100000",
                            698 => "111001100",
                            699 => "001000010",
                            700 => "010101110",
                            701 => "000010000",
                            702 => "000000000",
                            703 => "010001011",
                            704 => "000000000",
                            705 => "000000000",
                            706 => "010000010",
                            707 => "101001100",
                            708 => "101111110",
                            709 => "010000000",
                            710 => "000000000",
                            711 => "010100010",
                            712 => "000001100",
                            713 => "000110110",
                            714 => "100110000",
                            715 => "000111110",
                            716 => "000011010",
                            717 => "010010000",
                            718 => "000101100",
                            719 => "000010100",
                            720 => "110100010",
                            721 => "111101010",
                            722 => "011010110",
                            723 => "000000010",
                            724 => "101110110",
                            725 => "110011000",
                            726 => "000110110",
                            727 => "111110000",
                            728 => "101011010",
                            729 => "111011000",
                            730 => "011101010",
                            731 => "011111110",
                            732 => "011100100",
                            733 => "011011010",
                            734 => "101010000",
                            735 => "010100000",
                            736 => "000110000",
                            737 => "000000010",
                            738 => "101001100",
                            739 => "000001110",
                            740 => "011110100",
                            741 => "000000000",
                            742 => "000000000",
                            743 => "000101110",
                            744 => "000000110",
                            745 => "000000110",
                            746 => "000000000",
                            747 => "000101000",
                            748 => "111000000",
                            749 => "011011000",
                            750 => "101100110",
                            751 => "000011010",
                            752 => "110110000",
                            753 => "101001000",
                            754 => "101111000",
                            755 => "011000110",
                            756 => "110111000",
                            757 => "111111100",
                            758 => "001111110",
                            759 => "110011010",
                            760 => "001000110",
                            761 => "001101010",
                            762 => "000110100",
                            763 => "010011100",
                            764 => "110000010",
                            765 => "001110100",
                            766 => "110101110",
                            767 => "100111000",
                            768 => "101101100",
                            769 => "110100000",
                            770 => "000101110",
                            771 => "010010110",
                            772 => "000010010",
                            773 => "000000000",
                            774 => "001001110",
                            775 => "100100000",
                            776 => "111001100",
                            777 => "001000010",
                            778 => "010101110",
                            779 => "000010000",
                            780 => "000000000",
                            781 => "010001011",
                            782 => "000000000",
                            783 => "000000000",
                            784 => "010000010",
                            785 => "110100010",
                            786 => "101001000",
                            787 => "010000000",
                            788 => "000000000",
                            789 => "010100100",
                            790 => "000001100",
                            791 => "111011110",
                            792 => "101100100",
                            793 => "000111110",
                            794 => "000011010",
                            795 => "010010000",
                            796 => "000101100",
                            797 => "000010100",
                            798 => "110100010",
                            799 => "111101010",
                            800 => "011010110",
                            801 => "000000010",
                            802 => "101110110",
                            803 => "111001110",
                            804 => "001010100",
                            805 => "110100000",
                            806 => "001010110",
                            807 => "001010010",
                            808 => "100110010",
                            809 => "000011100",
                            810 => "101000100",
                            811 => "011110000",
                            812 => "111001110",
                            813 => "010100000",
                            814 => "000110000",
                            815 => "000001000",
                            816 => "010010100",
                            817 => "011110010",
                            818 => "110011110",
                            819 => "000000000",
                            820 => "000000000",
                            821 => "000101110",
                            822 => "000000110",
                            823 => "000000110",
                            824 => "000000000",
                            825 => "000101000",
                            826 => "111010100",
                            827 => "000111010",
                            828 => "001100100",
                            829 => "000000000",
                            830 => "111000110",
                            831 => "100101010",
                            832 => "111011100",
                            833 => "101101110",
                            834 => "001010100",
                            835 => "000101100",
                            836 => "111011010",
                            837 => "010100010",
                            838 => "001010110",
                            839 => "101001010",
                            840 => "111000100",
                            841 => "100000100",
                            842 => "000010110",
                            843 => "000101100",
                            844 => "111001000",
                            845 => "000000000",
                            846 => "000000000",
                            847 => "000011000",
                            848 => "100111110",
                            849 => "111100100",
                            850 => "010101110",
                            851 => "100111000",
                            852 => "101101100",
                            853 => "110100000",
                            854 => "000101110",
                            855 => "010010110",
                            856 => "000010010",
                            857 => "000010000",
                            858 => "000000000",
                            859 => "010001011",
                            860 => "000000000",
                            861 => "000000000",
                            862 => "001010000",
                            863 => "100101010",
                            864 => "001011010",
                            865 => "010000000",
                            866 => "000000000",
                            867 => "100000000",
                            868 => "000001100",
                            869 => "001110010",
                            870 => "110111000",
                            871 => "000010100",
                            872 => "110100010",
                            873 => "111101010",
                            874 => "011010110",
                            875 => "101000100",
                            876 => "100111110",
                            877 => "100010000",
                            878 => "111010100",
                            879 => "111001110",
                            880 => "000101110",
                            881 => "000000010",
                            882 => "101110110",
                            883 => "011101110",
                            884 => "001011010",
                            885 => "101000110",
                            886 => "110001100",
                            887 => "000011110",
                            888 => "001010110",
                            889 => "100010100",
                            890 => "000011000",
                            891 => "010100000",
                            892 => "000100000",
                            893 => "000000010",
                            894 => "111111100",
                            895 => "111001010",
                            896 => "000100010",
                            897 => "000000000",
                            898 => "000000000",
                            899 => "100111000",
                            900 => "101101100",
                            901 => "110100000",
                            902 => "000101110",
                            903 => "010010110",
                            904 => "000010010",
                            905 => "000000000",
                            906 => "001001110",
                            907 => "100100000",
                            908 => "111001100",
                            909 => "001000010",
                            910 => "010101110",
                            911 => "000010000",
                            912 => "000000000",
                            913 => "010001011",
                            914 => "000000000",
                            915 => "000000000",
                            916 => "010000010",
                            917 => "010011000",
                            918 => "000110110",
                            919 => "010000000",
                            920 => "000000000",
                            921 => "010100010",
                            922 => "000001100",
                            923 => "011101100",
                            924 => "001111000",
                            925 => "000111110",
                            926 => "000011010",
                            927 => "010010000",
                            928 => "000101100",
                            929 => "000010100",
                            930 => "110100010",
                            931 => "111101010",
                            932 => "011010110",
                            933 => "000000010",
                            934 => "101110110",
                            935 => "111001110",
                            936 => "001011000",
                            937 => "111110010",
                            938 => "001110000",
                            939 => "010000100",
                            940 => "100000100",
                            941 => "101000110",
                            942 => "011100100",
                            943 => "001000100",
                            944 => "001011110",
                            945 => "010100000",
                            946 => "000110000",
                            947 => "000000010",
                            948 => "001011000",
                            949 => "000010110",
                            950 => "001001110",
                            951 => "000000000",
                            952 => "000000000",
                            953 => "000101110",
                            954 => "000000110",
                            955 => "000000110",
                            956 => "000000000",
                            957 => "000101000",
                            958 => "111111000",
                            959 => "101101110",
                            960 => "101000000",
                            961 => "011110110",
                            962 => "010100100",
                            963 => "000000110",
                            964 => "101010100",
                            965 => "100110100",
                            966 => "110101100",
                            967 => "111111010",
                            968 => "001010110",
                            969 => "011101110",
                            970 => "010000110",
                            971 => "011010100",
                            972 => "010011000",
                            973 => "111110100",
                            974 => "111111010",
                            975 => "111000100",
                            976 => "100011100",
                            977 => "100111000",
                            978 => "101101100",
                            979 => "110100000",
                            980 => "000101110",
                            981 => "010010110",
                            982 => "000010010",
                            983 => "000000000",
                            984 => "001001110",
                            985 => "100100000",
                            986 => "111001100",
                            987 => "001000010",
                            988 => "010101110",
                            989 => "000010000",
                            990 => "000000000",
                            991 => "010001011",
                            992 => "000000000",
                            993 => "000000000",
                            994 => "010000010",
                            995 => "001001110",
                            996 => "101110110",
                            997 => "010000000",
                            998 => "000000000",
                            999 => "010100100",
                            1000 => "000001100",
                            1001 => "100110010",
                            1002 => "100111000",
                            1003 => "000111110",
                            1004 => "000011010",
                            1005 => "010010000",
                            1006 => "000101100",
                            1007 => "000010100",
                            1008 => "110100010",
                            1009 => "111101010",
                            1010 => "011010110",
                            1011 => "000000010",
                            1012 => "101110110",
                            1013 => "111001110",
                            1014 => "001010010",
                            1015 => "001001010",
                            1016 => "111000010",
                            1017 => "000111110",
                            1018 => "010010010",
                            1019 => "001100010",
                            1020 => "000010100",
                            1021 => "110001110",
                            1022 => "000000000",
                            1023 => "010100000",
                            1024 => "000110000",
                            1025 => "000000010",
                            1026 => "001001110",
                            1027 => "110100010",
                            1028 => "010000010",
                            1029 => "000000000",
                            1030 => "000000000",
                            1031 => "000101110",
                            1032 => "000000110",
                            1033 => "000000110",
                            1034 => "000000000",
                            1035 => "000101000",
                            1036 => "001111110",
                            1037 => "011101010",
                            1038 => "011010110",
                            1039 => "001111100",
                            1040 => "011101000",
                            1041 => "101010110",
                            1042 => "000000000",
                            1043 => "100111110",
                            1044 => "111101010",
                            1045 => "011110000",
                            1046 => "000000110",
                            1047 => "101100000",
                            1048 => "101001010",
                            1049 => "001111110",
                            1050 => "000101010",
                            1051 => "011110110",
                            1052 => "001101010",
                            1053 => "011000000",
                            1054 => "110001000",
                            1055 => "000000000",
                            1056 => "000000000",
                            1057 => "000011000",
                            1058 => "100111110",
                            1059 => "111100100",
                            1060 => "010101110",
                            1061 => "100111000",
                            1062 => "101101100",
                            1063 => "110100000",
                            1064 => "000101110",
                            1065 => "010010110",
                            1066 => "000010010",
                            1067 => "000010000",
                            1068 => "000000000",
                            1069 => "010001011",
                            1070 => "000000000",
                            1071 => "000000000",
                            1072 => "001010000",
                            1073 => "111100100",
                            1074 => "011010100",
                            1075 => "010000000",
                            1076 => "000000000",
                            1077 => "100000000",
                            1078 => "000001100",
                            1079 => "101000010",
                            1080 => "000001010",
                            1081 => "000010100",
                            1082 => "110100010",
                            1083 => "111101010",
                            1084 => "011010110",
                            1085 => "000111110",
                            1086 => "000011010",
                            1087 => "010010000",
                            1088 => "000101100",
                            1089 => "111001110",
                            1090 => "001011000",
                            1091 => "000000010",
                            1092 => "101110110",
                            1093 => "101000110",
                            1094 => "011100100",
                            1095 => "001000100",
                            1096 => "001011110",
                            1097 => "111110010",
                            1098 => "001110000",
                            1099 => "010000100",
                            1100 => "100110110",
                            1101 => "010100000",
                            1102 => "000100000",
                            1103 => "000000100",
                            1104 => "000000000",
                            1105 => "010111000",
                            1106 => "000101110",
                            1107 => "000000000",
                            1108 => "000000000",
                            1109 => "000000000",
                            1110 => "000000000",
                            1111 => "000011000",
                            1112 => "100111110",
                            1113 => "111100100",
                            1114 => "010101110",
                            1115 => "100111000",
                            1116 => "101101100",
                            1117 => "110100000",
                            1118 => "000101110",
                            1119 => "010010110",
                            1120 => "000010010",
                            1121 => "000010000",
                            1122 => "000000000",
                            1123 => "010001011",
                            1124 => "000000000",
                            1125 => "000000000",
                            1126 => "001010000",
                            1127 => "111100100",
                            1128 => "011011000",
                            1129 => "010000000",
                            1130 => "000000000",
                            1131 => "100000000",
                            1132 => "000001100",
                            1133 => "101000010",
                            1134 => "000000110",
                            1135 => "000010100",
                            1136 => "110100010",
                            1137 => "111101010",
                            1138 => "011010110",
                            1139 => "000111110",
                            1140 => "000011010",
                            1141 => "010010000",
                            1142 => "000101100",
                            1143 => "110011000",
                            1144 => "000110110",
                            1145 => "000000010",
                            1146 => "101110110",
                            1147 => "011111110",
                            1148 => "011100100",
                            1149 => "011011010",
                            1150 => "101010000",
                            1151 => "111110000",
                            1152 => "101011010",
                            1153 => "111011000",
                            1154 => "100011100",
                            1155 => "010100000",
                            1156 => "000100000",
                            1157 => "000000010",
                            1158 => "111111010",
                            1159 => "101001100",
                            1160 => "010010010",
                            1161 => "000000000",
                            1162 => "000000000",
                            1163 => "000000000",
                            1164 => "000000000",
                            1165 => "000011000",
                            1166 => "100111110",
                            1167 => "111100100",
                            1168 => "010101110",
                            1169 => "100111000",
                            1170 => "101101100",
                            1171 => "110100000",
                            1172 => "000101110",
                            1173 => "010010110",
                            1174 => "000010010",
                            1175 => "000010000",
                            1176 => "000000000",
                            1177 => "010001011",
                            1178 => "000000000",
                            1179 => "000000000",
                            1180 => "001010000",
                            1181 => "111100100",
                            1182 => "011010110",
                            1183 => "010000000",
                            1184 => "000000000",
                            1185 => "100000000",
                            1186 => "000001100",
                            1187 => "101000010",
                            1188 => "000001000",
                            1189 => "000010100",
                            1190 => "110100010",
                            1191 => "111101010",
                            1192 => "011010110",
                            1193 => "000111110",
                            1194 => "000011010",
                            1195 => "010010000",
                            1196 => "000101100",
                            1197 => "111001110",
                            1198 => "001010100",
                            1199 => "000000010",
                            1200 => "101110110",
                            1201 => "000011100",
                            1202 => "101000100",
                            1203 => "011110000",
                            1204 => "111001110",
                            1205 => "110100000",
                            1206 => "001010110",
                            1207 => "001010010",
                            1208 => "101100100",
                            1209 => "010100000",
                            1210 => "000100000",
                            1211 => "000000010",
                            1212 => "111111110",
                            1213 => "110111000",
                            1214 => "001010000",
                            1215 => "000000000",
                            1216 => "000000000",
                            1217 => "000000000",
                            1218 => "000000000",
                            1219 => "000011000",
                            1220 => "100111110",
                            1221 => "111100100",
                            1222 => "010101110",
                            1223 => "100111000",
                            1224 => "101101100",
                            1225 => "110100000",
                            1226 => "000101110",
                            1227 => "010010110",
                            1228 => "000010010",
                            1229 => "000010000",
                            1230 => "000000000",
                            1231 => "010001011",
                            1232 => "000000000",
                            1233 => "000000000",
                            1234 => "001010000",
                            1235 => "111100100",
                            1236 => "011011010",
                            1237 => "010000000",
                            1238 => "000000000",
                            1239 => "100000000",
                            1240 => "000001100",
                            1241 => "101000010",
                            1242 => "000000100",
                            1243 => "000010100",
                            1244 => "110100010",
                            1245 => "111101010",
                            1246 => "011010110",
                            1247 => "000111110",
                            1248 => "000011010",
                            1249 => "010010000",
                            1250 => "000101100",
                            1251 => "111001110",
                            1252 => "001010010",
                            1253 => "000000010",
                            1254 => "101110110",
                            1255 => "001100010",
                            1256 => "000010100",
                            1257 => "110001110",
                            1258 => "000000000",
                            1259 => "001001010",
                            1260 => "111000010",
                            1261 => "000111110",
                            1262 => "011000100",
                            1263 => "010100000",
                            1264 => "000100000",
                            1265 => "000000100",
                            1266 => "000000000",
                            1267 => "001000000",
                            1268 => "010000100",
                            1269 => "000000000",
                            1270 => "000000000",
                            1271 => "100111000",
                            1272 => "101101100",
                            1273 => "110100000",
                            1274 => "000101110",
                            1275 => "010010110",
                            1276 => "000010010",
                            1277 => "000000000",
                            1278 => "001001110",
                            1279 => "100100000",
                            1280 => "111001100",
                            1281 => "001000010",
                            1282 => "010101110",
                            1283 => "000010000",
                            1284 => "000000000",
                            1285 => "010001011",
                            1286 => "000000000",
                            1287 => "000000010",
                            1288 => "001000000",
                            1289 => "110111000",
                            1290 => "010010110",
                            1291 => "010000000",
                            1292 => "000000000",
                            1293 => "001101000",
                            1294 => "000001100",
                            1295 => "001111010",
                            1296 => "110001100",
                            1297 => "101000100",
                            1298 => "100111110",
                            1299 => "100010000",
                            1300 => "111010100",
                            1301 => "000010100",
                            1302 => "110100010",
                            1303 => "111101010",
                            1304 => "011010110",
                            1305 => "000000010",
                            1306 => "101110110",
                            1307 => "111001110",
                            1308 => "000101110",
                            1309 => "000011110",
                            1310 => "001010110",
                            1311 => "100010100",
                            1312 => "000011000",
                            1313 => "011101110",
                            1314 => "001011010",
                            1315 => "101000110",
                            1316 => "110001100",
                            1317 => "010100000",
                            1318 => "000110000",
                            1319 => "000000000",
                            1320 => "010101000",
                            1321 => "110011100",
                            1322 => "001100000",
                            1323 => "000000000",
                            1324 => "000000000",
                            1325 => "000101110",
                            1326 => "000000110",
                            1327 => "000000110",
                            1328 => "000000000",
                            1329 => "111100110",
                            1330 => "110001100",
                            1331 => "100101100",
                            1332 => "111110110",
                            1333 => "001111010",
                            1334 => "001000000",
                            1335 => "000011110",
                            1336 => "010010110",
                            1337 => "101000100",
                            1338 => "101101100",
                            1339 => "011001000",
                            1340 => "101111010",
                            1341 => "101101110",
                            1342 => "110110010",
                            1343 => "001011000",
                            1344 => "111100010",
                            1345 => "111110000",
                            1346 => "001001100",
                            1347 => "110000110",
                            1348 => "000011010",
                            1349 => "000001000",
                            1350 => "111000100",
                            1351 => "001111100",
                            1352 => "111111000",
                            1353 => "001011110",
                            1354 => "000100100",
                            1355 => "101110010",
                            1356 => "010101000",
                            1357 => "000110100",
                            1358 => "000101100",
                            1359 => "100010100",
                            1360 => "111101110",
                            1361 => "011001100",
                            1362 => "110100000",
                            1363 => "101111110",
                            1364 => "110110000",
                            1365 => "101110000",
                            1366 => "101010000",
                            1367 => "001001000",
                            1368 => "101010100",
                            1369 => "100100000",
                            1370 => "111101100",
                            1371 => "111010000",
                            1372 => "101110000",
                            1373 => "010110100",
                            1374 => "000011010",
                            1375 => "101110110",
                            1376 => "110000010",
                            1377 => "001110010",
                            1378 => "100000110",
                            1379 => "000111010",
                            1380 => "000010100",
                            1381 => "101000110",
                            1382 => "101000000",
                            1383 => "111000010",
                            1384 => "101110110",
                            1385 => "010101010",
                            1386 => "001100000",
                            1387 => "111001010",
                            1388 => "100100010",
                            1389 => "101110010",
                            1390 => "001110000",
                            1391 => "111101000",
                            1392 => "011011010",
                            1393 => "001011010",
                            1394 => "111101110",
                            1395 => "001110010",
                            1396 => "000111100",
                            1397 => "111101010",
                            1398 => "100010000",
                            1399 => "001011100",
                            1400 => "011111000",
                            1401 => "000000100",
                            1402 => "000111110",
                            1403 => "100010000",
                            1404 => "001011010",
                            1405 => "110001110",
                            1406 => "010011000",
                            1407 => "011110010",
                            1408 => "010111100",
                            1409 => "101000010",
                            1410 => "100111000",
                            1411 => "010011110",
                            1412 => "111000000",
                            1413 => "000010010",
                            1414 => "001100010",
                            1415 => "111100010",
                            1416 => "110001000",
                            1417 => "011100100",
                            1418 => "010110010",
                            1419 => "100101110",
                            1420 => "110110000",
                            1421 => "111011110",
                            1422 => "001010010",
                            1423 => "010100100",
                            1424 => "101011100",
                            1425 => "101010000",
                            1426 => "100001100",
                            1427 => "010100010",
                            1428 => "101000000",
                            1429 => "011011010",
                            1430 => "101000010",
                            1431 => "101001000",
                            1432 => "100100010",
                            1433 => "001011010",
                            1434 => "111101010",
                            1435 => "000110000",
                            1436 => "001011000",
                            1437 => "101010100",
                            1438 => "100010010",
                            1439 => "110010000",
                            1440 => "000111110",
                            1441 => "000110110",
                            1442 => "101111000",
                            1443 => "000101010",
                            1444 => "011101010",
                            1445 => "010001000",
                            1446 => "000110010",
                            1447 => "001101110",
                            1448 => "000000010",
                            1449 => "011001110",
                            1450 => "101110100",
                            1451 => "000110110",
                            1452 => "101101110",
                            1453 => "111011010",
                            1454 => "010111110",
                            1455 => "111101100",
                            1456 => "100111110",
                            1457 => "010111010",
                            1458 => "011010010",
                            1459 => "101001010",
                            1460 => "100100100",
                            1461 => "101101000",
                            1462 => "111110000",
                            1463 => "000110000",
                            1464 => "110010110",
                            1465 => "011011110",
                            1466 => "110001010",
                            1467 => "101000010",
                            1468 => "000000110",
                            1469 => "001001100",
                            1470 => "011110110",
                            1471 => "100111100",
                            1472 => "110111000",
                            1473 => "011111100",
                            1474 => "110000010",
                            1475 => "110000100",
                            1476 => "010011000",
                            1477 => "001010110",
                            1478 => "100010110",
                            1479 => "111100100",
                            1480 => "001111100",
                            1481 => "000011000",
                            1482 => "011010000",
                            1483 => "110100000",
                            1484 => "110001010",
                            1485 => "010001000",
                            1486 => "100100110",
                            1487 => "011100110",
                            1488 => "100110000",
                            1489 => "101010100",
                            1490 => "110000010",
                            1491 => "000010000",
                            1492 => "011001010",
                            1493 => "011010000",
                            1494 => "110000010",
                            1495 => "010001000",
                            1496 => "110001010",
                            1497 => "100010010",
                            1498 => "110010000",
                            1499 => "111000100",
                            1500 => "111101000",
                            1501 => "110001010",
                            1502 => "110101100",
                            1503 => "100111100",
                            1504 => "110110000",
                            1505 => "101001000",
                            1506 => "011010010",
                            1507 => "111000110",
                            1508 => "001101110",
                            1509 => "010001000",
                            1510 => "100101110",
                            1511 => "011001000",
                            1512 => "011000100",
                            1513 => "001101000",
                            1514 => "101011100",
                            1515 => "001001100",
                            1516 => "000101000",
                            1517 => "000100100",
                            1518 => "000100100",
                            1519 => "110101010",
                            1520 => "010111100",
                            1521 => "111000110",
                            1522 => "010011110",
                            1523 => "010001100",
                            1524 => "110000010",
                            1525 => "110000110",
                            1526 => "110110000",
                            1527 => "101001010",
                            1528 => "001010100",
                            1529 => "010110110",
                            1530 => "010001000",
                            1531 => "111011010",
                            1532 => "010001000",
                            1533 => "100001000",
                            1534 => "111100110",
                            1535 => "011001000",
                            1536 => "001011100",
                            1537 => "001010010",
                            1538 => "000100110",
                            1539 => "101000110",
                            1540 => "100011000",
                            1541 => "110010100",
                            1542 => "110011010",
                            1543 => "111000010",
                            1544 => "001000110",
                            1545 => "000000100",
                            1546 => "110001010",
                            1547 => "100111010",
                            1548 => "001010000",
                            1549 => "110100110",
                            1550 => "101111010",
                            1551 => "100001100",
                            1552 => "110100110",
                            1553 => "101011000",
                            1554 => "001010010",
                            1555 => "110110000",
                            1556 => "101101100",
                            1557 => "111011000",
                            1558 => "011100100",
                            1559 => "111110000",
                            1560 => "101100110",
                            1561 => "010110110",
                            1562 => "110011000",
                            1563 => "111001010",
                            1564 => "001110100",
                            1565 => "001001100",
                            1566 => "111000110",
                            1567 => "111000000",
                            1568 => "011101010",
                            1569 => "110000000",
                            1570 => "100011100",
                            1571 => "000000110",
                            1572 => "100100110",
                            1573 => "000000000",
                            1574 => "000000000",
                            1575 => "000011000",
                            1576 => "100111110",
                            1577 => "111100100",
                            1578 => "010101110",
                            1579 => "100111000",
                            1580 => "101101100",
                            1581 => "110100000",
                            1582 => "000101110",
                            1583 => "010010110",
                            1584 => "000010010",
                            1585 => "000010000",
                            1586 => "000000000",
                            1587 => "010001011",
                            1588 => "000000000",
                            1589 => "000000000",
                            1590 => "001010000",
                            1591 => "100101010",
                            1592 => "001011100",
                            1593 => "010000000",
                            1594 => "000000000",
                            1595 => "100000000",
                            1596 => "000001100",
                            1597 => "001110010",
                            1598 => "110110110",
                            1599 => "000010100",
                            1600 => "110100010",
                            1601 => "111101010",
                            1602 => "011010110",
                            1603 => "101000100",
                            1604 => "100111110",
                            1605 => "100010000",
                            1606 => "111010100",
                            1607 => "111001110",
                            1608 => "000101110",
                            1609 => "000000010",
                            1610 => "101110110",
                            1611 => "011101110",
                            1612 => "001011010",
                            1613 => "101000110",
                            1614 => "110001100",
                            1615 => "000011110",
                            1616 => "001010110",
                            1617 => "100010110",
                            1618 => "000001000",
                            1619 => "010100000",
                            1620 => "000100000",
                            1621 => "000000010",
                            1622 => "111111010",
                            1623 => "111001000",
                            1624 => "000110100",
                            1625 => "000000000",
                            1626 => "000000000",
                            1627 => "100111000",
                            1628 => "101101100",
                            1629 => "110100000",
                            1630 => "000101110",
                            1631 => "010010110",
                            1632 => "000010010",
                            1633 => "000000000",
                            1634 => "001001110",
                            1635 => "100100000",
                            1636 => "111001100",
                            1637 => "001000010",
                            1638 => "010101110",
                            1639 => "000010000",
                            1640 => "000000000",
                            1641 => "010001011",
                            1642 => "000000000",
                            1643 => "000000000",
                            1644 => "110100110",
                            1645 => "110111000",
                            1646 => "010011000",
                            1647 => "010000000",
                            1648 => "000000000",
                            1649 => "001101000",
                            1650 => "000001100",
                            1651 => "001111100",
                            1652 => "000100100",
                            1653 => "101000100",
                            1654 => "100111110",
                            1655 => "100010000",
                            1656 => "111010100",
                            1657 => "000010100",
                            1658 => "110100010",
                            1659 => "111101010",
                            1660 => "011010110",
                            1661 => "000000010",
                            1662 => "101110110",
                            1663 => "111001110",
                            1664 => "000101110",
                            1665 => "000011110",
                            1666 => "001010110",
                            1667 => "100010110",
                            1668 => "000001000",
                            1669 => "011101110",
                            1670 => "001011010",
                            1671 => "101000110",
                            1672 => "110001100",
                            1673 => "010100000",
                            1674 => "000110000",
                            1675 => "000000000",
                            1676 => "010101000",
                            1677 => "000101110",
                            1678 => "100101000",
                            1679 => "000000000",
                            1680 => "000000000",
                            1681 => "000101110",
                            1682 => "000000110",
                            1683 => "000000110",
                            1684 => "000000000",
                            1685 => "101001100",
                            1686 => "110001000",
                            1687 => "111000100",
                            1688 => "010110100",
                            1689 => "011010110",
                            1690 => "010011010",
                            1691 => "110000110",
                            1692 => "001111000",
                            1693 => "101111010",
                            1694 => "111000000",
                            1695 => "100111110",
                            1696 => "101000100",
                            1697 => "011100010",
                            1698 => "001001110",
                            1699 => "100010010",
                            1700 => "100101110",
                            1701 => "010111100",
                            1702 => "100000010",
                            1703 => "011001100",
                            1704 => "100110010",
                            1705 => "001011000",
                            1706 => "000000010",
                            1707 => "101110110",
                            1708 => "000100110",
                            1709 => "111000000",
                            1710 => "001100110",
                            1711 => "101100000",
                            1712 => "111011000",
                            1713 => "100101000",
                            1714 => "010111110",
                            1715 => "111101110",
                            1716 => "011000010",
                            1717 => "001111010",
                            1718 => "111000100",
                            1719 => "000011010",
                            1720 => "000100100",
                            1721 => "100111110",
                            1722 => "100001110",
                            1723 => "100100100",
                            1724 => "000101010",
                            1725 => "101111110",
                            1726 => "010100100",
                            1727 => "100011010",
                            1728 => "001111110",
                            1729 => "110011010",
                            1730 => "101010000",
                            1731 => "111000010",
                            1732 => "111111110",
                            1733 => "011001110",
                            1734 => "110100110",
                            1735 => "100001110",
                            1736 => "010110010",
                            1737 => "011000000",
                            1738 => "010010010",
                            1739 => "110011010",
                            1740 => "011010110",
                            1741 => "000011110",
                            1742 => "011000100",
                            1743 => "101110100",
                            1744 => "101101110",
                            1745 => "001100110",
                            1746 => "011010010",
                            1747 => "111101110",
                            1748 => "100001100",
                            1749 => "000010000",
                            1750 => "011010010",
                            1751 => "010011100",
                            1752 => "100001010",
                            1753 => "111000010",
                            1754 => "001001010",
                            1755 => "001111000",
                            1756 => "000100000",
                            1757 => "101110010",
                            1758 => "000011000",
                            1759 => "010111100",
                            1760 => "101110010",
                            1761 => "010111100",
                            1762 => "010000110",
                            1763 => "101001110",
                            1764 => "001001000",
                            1765 => "110000100",
                            1766 => "001011010",
                            1767 => "010111000",
                            1768 => "100100100",
                            1769 => "110100000",
                            1770 => "101010000",
                            1771 => "100000110",
                            1772 => "111111100",
                            1773 => "011100100",
                            1774 => "001011100",
                            1775 => "100111110",
                            1776 => "101010000",
                            1777 => "001101110",
                            1778 => "001001100",
                            1779 => "111001110",
                            1780 => "001111010",
                            1781 => "011011010",
                            1782 => "010010110",
                            1783 => "010000010",
                            1784 => "100010000",
                            1785 => "001011110",
                            1786 => "011011100",
                            1787 => "010001100",
                            1788 => "111100110",
                            1789 => "110110100",
                            1790 => "110010110",
                            1791 => "111011010",
                            1792 => "010000000",
                            1793 => "101010110",
                            1794 => "001100100",
                            1795 => "001110110",
                            1796 => "000001000",
                            1797 => "000111010",
                            1798 => "111001000",
                            1799 => "001100010",
                            1800 => "100101100",
                            1801 => "000101100",
                            1802 => "011000110",
                            1803 => "101111010",
                            1804 => "011101100",
                            1805 => "101111000",
                            1806 => "010101110",
                            1807 => "010011010",
                            1808 => "111100100",
                            1809 => "111111110",
                            1810 => "111110000",
                            1811 => "111010010",
                            1812 => "110101100",
                            1813 => "001110000",
                            1814 => "011110100",
                            1815 => "101110110",
                            1816 => "000000100",
                            1817 => "001011000",
                            1818 => "011001100",
                            1819 => "010100010",
                            1820 => "000100100",
                            1821 => "000111000",
                            1822 => "010101100",
                            1823 => "110010100",
                            1824 => "111101000",
                            1825 => "101101010",
                            1826 => "001001000",
                            1827 => "000010010",
                            1828 => "100101010",
                            1829 => "010010100",
                            1830 => "101001110",
                            1831 => "101010100",
                            1832 => "010110010",
                            1833 => "110000000",
                            1834 => "000000000",
                            1835 => "011001010",
                            1836 => "110011010",
                            1837 => "101011110",
                            1838 => "000101000",
                            1839 => "110101010",
                            1840 => "001100010",
                            1841 => "101110110",
                            1842 => "101011010",
                            1843 => "000011100",
                            1844 => "110100010",
                            1845 => "110001100",
                            1846 => "101110010",
                            1847 => "000100000",
                            1848 => "000001000",
                            1849 => "010110000",
                            1850 => "100110100",
                            1851 => "100000000",
                            1852 => "000000000",
                            1853 => "000000000",
                            1854 => "000011000",
                            1855 => "100111110",
                            1856 => "111100100",
                            1857 => "010101110",
                            1858 => "100111000",
                            1859 => "101101100",
                            1860 => "110100000",
                            1861 => "000101110",
                            1862 => "010010110",
                            1863 => "000010010",
                            1864 => "000010000",
                            1865 => "000000000",
                            1866 => "010001011",
                            1867 => "000000000",
                            1868 => "000000000",
                            1869 => "001010000",
                            1870 => "100101010",
                            1871 => "001011110",
                            1872 => "010000000",
                            1873 => "000000000",
                            1874 => "100000000",
                            1875 => "000001100",
                            1876 => "001110010",
                            1877 => "110110100",
                            1878 => "000010100",
                            1879 => "110100010",
                            1880 => "111101010",
                            1881 => "011010110",
                            1882 => "101000100",
                            1883 => "100111110",
                            1884 => "100010000",
                            1885 => "111010100",
                            1886 => "111001110",
                            1887 => "000101110",
                            1888 => "000000010",
                            1889 => "101110110",
                            1890 => "011101110",
                            1891 => "001011010",
                            1892 => "101000110",
                            1893 => "110001100",
                            1894 => "000011110",
                            1895 => "001010110",
                            1896 => "100010110",
                            1897 => "101011110",
                            1898 => "010100000",
                            1899 => "000100000",
                            1900 => "000000010",
                            1901 => "111111000",
                            1902 => "111000110",
                            1903 => "011100000",
                            1904 => "000000000",
                            1905 => "000000000",
                            1906 => "000000000",
                            1907 => "000000000",
                            1908 => "000011000",
                            1909 => "100111110",
                            1910 => "111100100",
                            1911 => "010101110",
                            1912 => "100111000",
                            1913 => "101101100",
                            1914 => "110100000",
                            1915 => "000101110",
                            1916 => "010010110",
                            1917 => "000010010",
                            1918 => "000010000",
                            1919 => "000000000",
                            1920 => "010001011",
                            1921 => "100110000",
                            1922 => "000000000",
                            1923 => "010001010",
                            1924 => "111100100",
                            1925 => "011011100",
                            1926 => "010000000",
                            1927 => "000000000",
                            1928 => "100000000",
                            1929 => "000001100",
                            1930 => "101000000",
                            1931 => "010011000",
                            1932 => "000010100",
                            1933 => "110100010",
                            1934 => "111101010",
                            1935 => "011010110",
                            1936 => "000111110",
                            1937 => "000011010",
                            1938 => "010010000",
                            1939 => "000101100",
                            1940 => "110011000",
                            1941 => "001100110",
                            1942 => "000000010",
                            1943 => "101110110",
                            1944 => "101000000",
                            1945 => "110101110",
                            1946 => "100100000",
                            1947 => "110000000",
                            1948 => "010010110",
                            1949 => "010101010",
                            1950 => "000101000",
                            1951 => "100001110",
                            1952 => "010100000",
                            1953 => "000110000",
                            1954 => "000000010",
                            1955 => "111111100",
                            1956 => "010001100",
                            1957 => "010010000",
                            1958 => "000000000",
                            1959 => "000000000",
                            1960 => "000101110",
                            1961 => "000000110",
                            1962 => "000000110",
                            1963 => "000000000",
                            1964 => "000110000",
                            1965 => "000101010",
                            1966 => "010100010",
                            1967 => "111001000",
                            1968 => "111110000",
                            1969 => "010111100",
                            1970 => "001110100",
                            1971 => "110010110",
                            1972 => "101110110",
                            1973 => "011011000",
                            1974 => "011010100",
                            1975 => "101101110",
                            1976 => "011100110",
                            1977 => "111110110",
                            1978 => "100011000",
                            1979 => "010110100",
                            1980 => "100001010",
                            1981 => "010011110",
                            1982 => "000111110",
                            1983 => "000100000",
                            1984 => "010011110",
                            1985 => "010010110",
                            1986 => "110110010",
                            1987 => "010110010",
                            1988 => "111101100",
                            1989 => "100111000",
                            1990 => "101101100",
                            1991 => "110100000",
                            1992 => "000101110",
                            1993 => "010010110",
                            1994 => "000010010",
                            1995 => "000000000",
                            1996 => "001001110",
                            1997 => "100100000",
                            1998 => "111001100",
                            1999 => "001000010",
                            2000 => "010101110",
                            2001 => "000010000",
                            2002 => "000000000",
                            2003 => "010001011",
                            2004 => "000000000",
                            2005 => "000000010",
                            2006 => "000111110",
                            2007 => "110111000",
                            2008 => "010011010",
                            2009 => "010000000",
                            2010 => "000000000",
                            2011 => "001101000",
                            2012 => "000001100",
                            2013 => "001111010",
                            2014 => "110001010",
                            2015 => "101000100",
                            2016 => "100111110",
                            2017 => "100010000",
                            2018 => "111010100",
                            2019 => "000010100",
                            2020 => "110100010",
                            2021 => "111101010",
                            2022 => "011010110",
                            2023 => "000000010",
                            2024 => "101110110",
                            2025 => "111001110",
                            2026 => "000101110",
                            2027 => "000011110",
                            2028 => "001010110",
                            2029 => "100010110",
                            2030 => "101011110",
                            2031 => "011101110",
                            2032 => "001011010",
                            2033 => "101000110",
                            2034 => "110001100",
                            2035 => "010100000",
                            2036 => "000110000",
                            2037 => "000000000",
                            2038 => "010101000",
                            2039 => "000100100",
                            2040 => "001010100",
                            2041 => "000000000",
                            2042 => "000000000",
                            2043 => "000101110",
                            2044 => "000000110",
                            2045 => "000000110",
                            2046 => "000000000",
                            2047 => "111100100",
                            2048 => "110110010",
                            2049 => "100110100",
                            2050 => "011110100",
                            2051 => "110000100",
                            2052 => "000010000",
                            2053 => "111011000",
                            2054 => "001100100",
                            2055 => "111001000",
                            2056 => "101100100",
                            2057 => "001100110",
                            2058 => "101010100",
                            2059 => "010010110",
                            2060 => "011001010",
                            2061 => "000001000",
                            2062 => "100011100",
                            2063 => "100111000",
                            2064 => "101010010",
                            2065 => "001010000",
                            2066 => "001101000",
                            2067 => "100010010",
                            2068 => "010011010",
                            2069 => "111110010",
                            2070 => "010011100",
                            2071 => "001111010",
                            2072 => "000010100",
                            2073 => "111011110",
                            2074 => "000110010",
                            2075 => "110010110",
                            2076 => "110110000",
                            2077 => "011110100",
                            2078 => "010111100",
                            2079 => "010101110",
                            2080 => "100111110",
                            2081 => "110101110",
                            2082 => "010000000",
                            2083 => "110110000",
                            2084 => "110000010",
                            2085 => "100100110",
                            2086 => "010100100",
                            2087 => "001010000",
                            2088 => "000100100",
                            2089 => "011110100",
                            2090 => "100110010",
                            2091 => "110011000",
                            2092 => "001100110",
                            2093 => "100001010",
                            2094 => "101010010",
                            2095 => "000010000",
                            2096 => "111111110",
                            2097 => "110011010",
                            2098 => "110111000",
                            2099 => "110011100",
                            2100 => "001001000",
                            2101 => "000000110",
                            2102 => "011111010",
                            2103 => "011000100",
                            2104 => "000010100",
                            2105 => "100110100",
                            2106 => "001001100",
                            2107 => "100111000",
                            2108 => "010011110",
                            2109 => "011001000",
                            2110 => "010101000",
                            2111 => "110001100",
                            2112 => "111110000",
                            2113 => "000101100",
                            2114 => "011001010",
                            2115 => "111101110",
                            2116 => "000011100",
                            2117 => "011010100",
                            2118 => "000000110",
                            2119 => "110000100",
                            2120 => "000100110",
                            2121 => "000011110",
                            2122 => "100010010",
                            2123 => "000010010",
                            2124 => "010001110",
                            2125 => "000101000",
                            2126 => "001000100",
                            2127 => "001100110",
                            2128 => "011111100",
                            2129 => "001101110",
                            2130 => "001010000",
                            2131 => "110001010",
                            2132 => "100000110",
                            2133 => "110101010",
                            2134 => "101110010",
                            2135 => "110101000",
                            2136 => "110101110",
                            2137 => "000011100",
                            2138 => "001110110",
                            2139 => "101000000",
                            2140 => "011011000",
                            2141 => "001110000",
                            2142 => "011111000",
                            2143 => "010111110",
                            2144 => "010001010",
                            2145 => "101100110",
                            2146 => "111111010",
                            2147 => "010100110",
                            2148 => "101001110",
                            2149 => "000110000",
                            2150 => "000001010",
                            2151 => "000011010",
                            2152 => "001100100",
                            2153 => "100111110",
                            2154 => "010111000",
                            2155 => "001001000",
                            2156 => "101111010",
                            2157 => "101010100",
                            2158 => "010111000",
                            2159 => "010110000",
                            2160 => "101000000",
                            2161 => "001000010",
                            2162 => "110100010",
                            2163 => "110001100",
                            2164 => "100100110",
                            2165 => "101000100",
                            2166 => "100101000",
                            2167 => "100101010",
                            2168 => "001010110",
                            2169 => "010101000",
                            2170 => "010001100",
                            2171 => "111101100",
                            2172 => "011011100",
                            2173 => "110011000",
                            2174 => "111001000",
                            2175 => "010011100",
                            2176 => "000101110",
                            2177 => "100011110",
                            2178 => "011101110",
                            2179 => "010010110",
                            2180 => "010001110",
                            2181 => "001110110",
                            2182 => "101001110",
                            2183 => "000100000",
                            2184 => "011111110",
                            2185 => "100000010",
                            2186 => "110100110",
                            2187 => "011001110",
                            2188 => "111101100",
                            2189 => "110001110",
                            2190 => "000010010",
                            2191 => "001001110",
                            2192 => "001000110",
                            2193 => "110001110",
                            2194 => "000100000",
                            2195 => "101011000",
                            2196 => "110010010",
                            2197 => "001111110",
                            2198 => "011111110",
                            2199 => "000001010",
                            2200 => "000011110",
                            2201 => "110000100",
                            2202 => "011000110",
                            2203 => "100100100",
                            2204 => "111100100",
                            2205 => "010100110",
                            2206 => "000000010",
                            2207 => "111000000",
                            2208 => "111101000",
                            2209 => "100010010",
                            2210 => "000011000",
                            2211 => "101010110",
                            2212 => "110100110",
                            2213 => "101011000",
                            2214 => "110100000",
                            2215 => "000111000",
                            2216 => "111100100",
                            2217 => "001001100",
                            2218 => "011100100",
                            2219 => "010011100",
                            2220 => "100010010",
                            2221 => "001101110",
                            2222 => "000000100",
                            2223 => "110110010",
                            2224 => "100010000",
                            2225 => "110100000",
                            2226 => "110001010",
                            2227 => "010001100",
                            2228 => "000100100",
                            2229 => "110010010",
                            2230 => "010010100",
                            2231 => "100101000",
                            2232 => "100011110",
                            2233 => "001110010",
                            2234 => "001001010",
                            2235 => "100010010",
                            2236 => "001101010",
                            2237 => "010010110",
                            2238 => "001111000",
                            2239 => "110101010",
                            2240 => "100010110",
                            2241 => "011011110",
                            2242 => "000111000",
                            2243 => "000101010",
                            2244 => "100010100",
                            2245 => "111000110",
                            2246 => "011001010",
                            2247 => "010000010",
                            2248 => "000101110",
                            2249 => "001100110",
                            2250 => "101000010",
                            2251 => "001101110",
                            2252 => "010101100",
                            2253 => "010111110",
                            2254 => "000110000",
                            2255 => "000111100",
                            2256 => "110101010",
                            2257 => "001100000",
                            2258 => "001110100",
                            2259 => "011101100",
                            2260 => "111001010",
                            2261 => "001010000",
                            2262 => "010111100",
                            2263 => "101111010",
                            2264 => "010100110",
                            2265 => "110110010",
                            2266 => "011001110",
                            2267 => "000111100",
                            2268 => "101010100",
                            2269 => "010000110",
                            2270 => "011001000",
                            2271 => "000000000",
                            2272 => "110101010",
                            2273 => "001010000",
                            2274 => "000100110",
                            2275 => "010011000",
                            2276 => "111010000",
                            2277 => "010101110",
                            2278 => "000110100",
                            2279 => "000001000",
                            2280 => "110111000",
                            2281 => "101000100",
                            2282 => "011011100",
                            2283 => "010111010",
                            2284 => "001011110",
                            2285 => "000011010",
                            2286 => "111101100",
                            2287 => "000101110",
                            2288 => "110001010",
                            2289 => "111011110",
                            2290 => "100111000",
                            2291 => "101101100",
                            2292 => "110100000",
                            2293 => "000101110",
                            2294 => "010010110",
                            2295 => "000010010",
                            2296 => "000000000",
                            2297 => "001001110",
                            2298 => "100100000",
                            2299 => "111001100",
                            2300 => "001000010",
                            2301 => "010101110",
                            2302 => "000010000",
                            2303 => "000000000",
                            2304 => "010001011",
                            2305 => "000000000",
                            2306 => "000000000",
                            2307 => "001010000",
                            2308 => "110001110",
                            2309 => "000011010",
                            2310 => "010000000",
                            2311 => "000000000",
                            2312 => "010100010",
                            2313 => "000001100",
                            2314 => "111110110",
                            2315 => "011000100",
                            2316 => "000111110",
                            2317 => "000011010",
                            2318 => "010010000",
                            2319 => "000101100",
                            2320 => "000010100",
                            2321 => "110100010",
                            2322 => "111101010",
                            2323 => "011010110",
                            2324 => "000000010",
                            2325 => "101110110",
                            2326 => "110011000",
                            2327 => "001100110",
                            2328 => "010010110",
                            2329 => "010101010",
                            2330 => "000101000",
                            2331 => "100001110",
                            2332 => "101000000",
                            2333 => "110101110",
                            2334 => "100100000",
                            2335 => "110111010",
                            2336 => "010100000",
                            2337 => "000100000",
                            2338 => "000000010",
                            2339 => "001001110",
                            2340 => "111001110",
                            2341 => "110011010",
                            2342 => "000000000",
                            2343 => "000000000",
                            2344 => "000000000",
                            2345 => "000000000",
                            2346 => "000011000",
                            2347 => "100111110",
                            2348 => "111100100",
                            2349 => "010101110",
                            2350 => "100111000",
                            2351 => "101101100",
                            2352 => "110100000",
                            2353 => "000101110",
                            2354 => "010010110",
                            2355 => "000010010",
                            2356 => "000010000",
                            2357 => "000000000",
                            2358 => "010001011",
                            2359 => "000000000",
                            2360 => "000000000",
                            2361 => "001010000",
                            2362 => "100101010",
                            2363 => "001100000",
                            2364 => "010000000",
                            2365 => "000000000",
                            2366 => "100000000",
                            2367 => "000001100",
                            2368 => "001110010",
                            2369 => "110110010",
                            2370 => "000010100",
                            2371 => "110100010",
                            2372 => "111101010",
                            2373 => "011010110",
                            2374 => "101000100",
                            2375 => "100111110",
                            2376 => "100010000",
                            2377 => "111010100",
                            2378 => "111001110",
                            2379 => "000101110",
                            2380 => "000000010",
                            2381 => "101110110",
                            2382 => "011101110",
                            2383 => "001011010",
                            2384 => "101000110",
                            2385 => "110001100",
                            2386 => "000011110",
                            2387 => "001010110",
                            2388 => "100011000",
                            2389 => "101001100",
                            2390 => "010100000",
                            2391 => "000100000",
                            2392 => "000000010",
                            2393 => "111111000",
                            2394 => "111000100",
                            2395 => "011110010",
                            2396 => "000000000",
                            2397 => "000000000",
                            2398 => "100111000",
                            2399 => "101101100",
                            2400 => "110100000",
                            2401 => "000101110",
                            2402 => "010010110",
                            2403 => "000010010",
                            2404 => "000000000",
                            2405 => "001001110",
                            2406 => "100100000",
                            2407 => "111001100",
                            2408 => "001000010",
                            2409 => "010101110",
                            2410 => "000010000",
                            2411 => "000000000",
                            2412 => "010001011",
                            2413 => "000000000",
                            2414 => "000000000",
                            2415 => "010000010",
                            2416 => "110001110",
                            2417 => "000011100",
                            2418 => "010000000",
                            2419 => "000000000",
                            2420 => "010100010",
                            2421 => "000001100",
                            2422 => "111110110",
                            2423 => "010010000",
                            2424 => "000111110",
                            2425 => "000011010",
                            2426 => "010010000",
                            2427 => "000101100",
                            2428 => "000010100",
                            2429 => "110100010",
                            2430 => "111101010",
                            2431 => "011010110",
                            2432 => "000000010",
                            2433 => "101110110",
                            2434 => "110011000",
                            2435 => "001100110",
                            2436 => "010010110",
                            2437 => "010101010",
                            2438 => "000101000",
                            2439 => "100001110",
                            2440 => "101000000",
                            2441 => "110101110",
                            2442 => "100100000",
                            2443 => "110111010",
                            2444 => "010100000",
                            2445 => "000110000",
                            2446 => "000000010",
                            2447 => "001001110",
                            2448 => "101100110",
                            2449 => "010001110",
                            2450 => "000000000",
                            2451 => "000000000",
                            2452 => "000101110",
                            2453 => "000000110",
                            2454 => "000000110",
                            2455 => "000000000",
                            2456 => "000101000",
                            2457 => "110110100",
                            2458 => "101011010",
                            2459 => "100110010",
                            2460 => "111010100",
                            2461 => "010000110",
                            2462 => "000101000",
                            2463 => "100010110",
                            2464 => "110000110",
                            2465 => "001100000",
                            2466 => "010101000",
                            2467 => "101000010",
                            2468 => "001110010",
                            2469 => "100001010",
                            2470 => "001011000",
                            2471 => "010110100",
                            2472 => "001001100",
                            2473 => "000101010",
                            2474 => "111100000",
                            2475 => "010101110",
                            2476 => "000000000",
                            2477 => "000000000",
                            2478 => "000011000",
                            2479 => "100111110",
                            2480 => "111100100",
                            2481 => "010101110",
                            2482 => "100111000",
                            2483 => "101101100",
                            2484 => "110100000",
                            2485 => "000101110",
                            2486 => "010010110",
                            2487 => "000010010",
                            2488 => "000010000",
                            2489 => "000000000",
                            2490 => "010001011",
                            2491 => "000000000",
                            2492 => "000000000",
                            2493 => "001010000",
                            2494 => "111100100",
                            2495 => "011011110",
                            2496 => "010000000",
                            2497 => "000000000",
                            2498 => "100000000",
                            2499 => "000001100",
                            2500 => "101000010",
                            2501 => "000000000",
                            2502 => "000010100",
                            2503 => "110100010",
                            2504 => "111101010",
                            2505 => "011010110",
                            2506 => "000111110",
                            2507 => "000011010",
                            2508 => "010010000",
                            2509 => "000101100",
                            2510 => "110011000",
                            2511 => "001100110",
                            2512 => "000000010",
                            2513 => "101110110",
                            2514 => "101000000",
                            2515 => "110101110",
                            2516 => "100100000",
                            2517 => "110111010",
                            2518 => "010010110",
                            2519 => "010101010",
                            2520 => "000101000",
                            2521 => "101000000",
                            2522 => "010100000",
                            2523 => "000100000",
                            2524 => "000000010",
                            2525 => "111111100",
                            2526 => "111001100",
                            2527 => "110111010",
                            2528 => "000000000",
                            2529 => "000000000",
                            2530 => "100111000",
                            2531 => "101101100",
                            2532 => "110100000",
                            2533 => "000101110",
                            2534 => "010010110",
                            2535 => "000010010",
                            2536 => "000000000",
                            2537 => "001001110",
                            2538 => "100100000",
                            2539 => "111001100",
                            2540 => "001000010",
                            2541 => "010101110",
                            2542 => "000010000",
                            2543 => "000000000",
                            2544 => "010001011",
                            2545 => "000000000",
                            2546 => "000000010",
                            2547 => "010011100",
                            2548 => "110111000",
                            2549 => "010011100",
                            2550 => "010000000",
                            2551 => "000000000",
                            2552 => "001101000",
                            2553 => "000001100",
                            2554 => "001111010",
                            2555 => "100101010",
                            2556 => "101000100",
                            2557 => "100111110",
                            2558 => "100010000",
                            2559 => "111010100",
                            2560 => "000010100",
                            2561 => "110100010",
                            2562 => "111101010",
                            2563 => "011010110",
                            2564 => "000000010",
                            2565 => "101110110",
                            2566 => "111001110",
                            2567 => "000101110",
                            2568 => "000011110",
                            2569 => "001010110",
                            2570 => "100011000",
                            2571 => "101001100",
                            2572 => "011101110",
                            2573 => "001011010",
                            2574 => "101000110",
                            2575 => "110001100",
                            2576 => "010100000",
                            2577 => "000110000",
                            2578 => "000000000",
                            2579 => "010101000",
                            2580 => "100110110",
                            2581 => "011110110",
                            2582 => "000000000",
                            2583 => "000000000",
                            2584 => "000101110",
                            2585 => "000000110",
                            2586 => "000000110",
                            2587 => "000000010",
                            2588 => "001000010",
                            2589 => "101101110",
                            2590 => "111101100",
                            2591 => "011000100",
                            2592 => "001100100",
                            2593 => "001011100",
                            2594 => "011010000",
                            2595 => "100111010",
                            2596 => "010110110",
                            2597 => "100011100",
                            2598 => "011010110",
                            2599 => "111111010",
                            2600 => "111001100",
                            2601 => "010000110",
                            2602 => "100011110",
                            2603 => "100110100",
                            2604 => "000101000",
                            2605 => "010111010",
                            2606 => "000110010",
                            2607 => "111010110",
                            2608 => "010110000",
                            2609 => "011110100",
                            2610 => "101001010",
                            2611 => "101000110",
                            2612 => "000111000",
                            2613 => "100110010",
                            2614 => "011111110",
                            2615 => "001110000",
                            2616 => "101001100",
                            2617 => "111000110",
                            2618 => "000011010",
                            2619 => "101100100",
                            2620 => "000001000",
                            2621 => "101110110",
                            2622 => "111010100",
                            2623 => "111011000",
                            2624 => "111100000",
                            2625 => "101000000",
                            2626 => "000100010",
                            2627 => "101100000",
                            2628 => "110110010",
                            2629 => "110100100",
                            2630 => "010010100",
                            2631 => "101101010",
                            2632 => "010011100",
                            2633 => "111000100",
                            2634 => "111111010",
                            2635 => "000110100",
                            2636 => "011010000",
                            2637 => "111101000",
                            2638 => "011000000",
                            2639 => "010011000",
                            2640 => "100011000",
                            2641 => "001010010",
                            2642 => "101000110",
                            2643 => "011011000",
                            2644 => "100100100",
                            2645 => "110000010",
                            2646 => "101110110",
                            2647 => "011001010",
                            2648 => "001011110",
                            2649 => "010111010",
                            2650 => "100110000",
                            2651 => "111001110",
                            2652 => "101010100",
                            2653 => "111011100",
                            2654 => "001111000",
                            2655 => "010101010",
                            2656 => "010000000",
                            2657 => "100100110",
                            2658 => "000110000",
                            2659 => "001110110",
                            2660 => "111011010",
                            2661 => "010100000",
                            2662 => "110011010",
                            2663 => "111111000",
                            2664 => "001010100",
                            2665 => "101111110",
                            2666 => "111011110",
                            2667 => "101100010",
                            2668 => "111010000",
                            2669 => "010111110",
                            2670 => "100001110",
                            2671 => "001111010",
                            2672 => "010010010",
                            2673 => "001101110",
                            2674 => "111011110",
                            2675 => "000100000",
                            2676 => "001000010",
                            2677 => "010110100",
                            2678 => "000010010",
                            2679 => "100001000",
                            2680 => "100000100",
                            2681 => "100100110",
                            2682 => "000111000",
                            2683 => "110010100",
                            2684 => "110101100",
                            2685 => "100000000",
                            2686 => "001010110",
                            2687 => "010101000",
                            2688 => "011011110",
                            2689 => "110110100",
                            2690 => "100101010",
                            2691 => "010100100",
                            2692 => "111011110",
                            2693 => "111001010",
                            2694 => "001110110",
                            2695 => "011011110",
                            2696 => "001001000",
                            2697 => "100011000",
                            2698 => "011111110",
                            2699 => "001001010",
                            2700 => "010011100",
                            2701 => "011010100",
                            2702 => "011110010",
                            2703 => "011010010",
                            2704 => "110111110",
                            2705 => "010111110",
                            2706 => "111000010",
                            2707 => "100110110",
                            2708 => "000111110",
                            2709 => "000000000",
                            2710 => "100110000",
                            2711 => "000110000",
                            2712 => "010111110",
                            2713 => "100010110",
                            2714 => "001110000",
                            2715 => "101011000",
                            2716 => "110001000",
                            2717 => "101101010",
                            2718 => "100101100",
                            2719 => "101110110",
                            2720 => "100111000",
                            2721 => "111110010",
                            2722 => "111011100",
                            2723 => "011110000",
                            2724 => "001111010",
                            2725 => "111010010",
                            2726 => "000110110",
                            2727 => "010101110",
                            2728 => "001010110",
                            2729 => "010110000",
                            2730 => "000100110",
                            2731 => "011111110",
                            2732 => "010011000",
                            2733 => "000001100",
                            2734 => "000011010",
                            2735 => "110000010",
                            2736 => "011010000",
                            2737 => "100000110",
                            2738 => "011111110",
                            2739 => "001101010",
                            2740 => "100101010",
                            2741 => "010010010",
                            2742 => "100101000",
                            2743 => "110010100",
                            2744 => "101011010",
                            2745 => "000010010",
                            2746 => "100111110",
                            2747 => "111010000",
                            2748 => "000011010",
                            2749 => "010010100",
                            2750 => "100000100",
                            2751 => "101010000",
                            2752 => "100100110",
                            2753 => "001110000",
                            2754 => "101000010",
                            2755 => "101100010",
                            2756 => "111011110",
                            2757 => "000001010",
                            2758 => "001100000",
                            2759 => "111010100",
                            2760 => "111100110",
                            2761 => "111010100",
                            2762 => "001101110",
                            2763 => "110111100",
                            2764 => "011000010",
                            2765 => "011001000",
                            2766 => "111000010",
                            2767 => "001111100",
                            2768 => "000100000",
                            2769 => "010011010",
                            2770 => "101000000",
                            2771 => "011001110",
                            2772 => "000101010",
                            2773 => "101000110",
                            2774 => "101011110",
                            2775 => "100101110",
                            2776 => "101110010",
                            2777 => "100100000",
                            2778 => "001001000",
                            2779 => "010010000",
                            2780 => "000011110",
                            2781 => "101100010",
                            2782 => "001101100",
                            2783 => "111101100",
                            2784 => "100001100",
                            2785 => "011010000",
                            2786 => "001000110",
                            2787 => "000010110",
                            2788 => "010100010",
                            2789 => "100000010",
                            2790 => "011111010",
                            2791 => "010110100",
                            2792 => "000010100",
                            2793 => "101111000",
                            2794 => "111001010",
                            2795 => "101011110",
                            2796 => "010100100",
                            2797 => "110100000",
                            2798 => "000110100",
                            2799 => "010101110",
                            2800 => "001110000",
                            2801 => "101000100",
                            2802 => "010111100",
                            2803 => "100110010",
                            2804 => "011000000",
                            2805 => "010000100",
                            2806 => "001010000",
                            2807 => "001010010",
                            2808 => "111100110",
                            2809 => "110110010",
                            2810 => "101000100",
                            2811 => "101100110",
                            2812 => "111111110",
                            2813 => "111001000",
                            2814 => "111101000",
                            2815 => "010001100",
                            2816 => "101100110",
                            2817 => "010111110",
                            2818 => "111111110",
                            2819 => "111010110",
                            2820 => "000000100",
                            2821 => "110110110",
                            2822 => "011010100",
                            2823 => "000110100",
                            2824 => "001100110",
                            2825 => "101010100",
                            2826 => "000001000",
                            2827 => "100000110",
                            2828 => "011101100",
                            2829 => "011111000",
                            2830 => "101101100",
                            2831 => "010001010",
                            2832 => "101101100",
                            2833 => "100100010",
                            2834 => "101101010",
                            2835 => "100011110",
                            2836 => "010000000",
                            2837 => "111001000",
                            2838 => "110110000",
                            2839 => "001000110",
                            2840 => "010101000",
                            2841 => "011110110",
                            2842 => "110011110",
                            2843 => "100111110",
                            2844 => "111010100",
                            2845 => "011010100",
                            2846 => "110110010",
                            2847 => "010011010",
                            2848 => "010011000",
                            2849 => "100000000",
                            2850 => "101101100",
                            2851 => "111001100",
                            2852 => "111111010",
                            2853 => "000100010",
                            2854 => "110101100",
                            2855 => "001110100",
                            2856 => "010110110",
                            2857 => "111111010",
                            2858 => "110001100",
                            2859 => "110011000",
                            2860 => "111101100",
                            2861 => "101001010",
                            2862 => "011001100",
                            2863 => "001110110",
                            2864 => "010110110",
                            2865 => "111110110",
                            2866 => "010111010",
                            2867 => "100101000",
                            2868 => "000010100",
                            2869 => "110011110",
                            2870 => "000101110",
                            2871 => "101001100",
                            2872 => "100110010",
                            2873 => "000010010",
                            2874 => "001010110",
                            2875 => "011011100",
                            2876 => "100010100",
                            2877 => "000000010",
                            2878 => "000000000",
                            2879 => "000000000",
                            2880 => "000011000",
                            2881 => "100111110",
                            2882 => "111100100",
                            2883 => "010101110",
                            2884 => "100111000",
                            2885 => "101101100",
                            2886 => "110100000",
                            2887 => "000101110",
                            2888 => "010010110",
                            2889 => "000010010",
                            2890 => "000010000",
                            2891 => "000000000",
                            2892 => "010001011",
                            2893 => "000000000",
                            2894 => "000000000",
                            2895 => "001010000",
                            2896 => "100101010",
                            2897 => "001100010",
                            2898 => "010000000",
                            2899 => "000000000",
                            2900 => "100000000",
                            2901 => "000001100",
                            2902 => "001110010",
                            2903 => "110110000",
                            2904 => "000010100",
                            2905 => "110100010",
                            2906 => "111101010",
                            2907 => "011010110",
                            2908 => "101000100",
                            2909 => "100111110",
                            2910 => "100010000",
                            2911 => "111010100",
                            2912 => "111001110",
                            2913 => "000101110",
                            2914 => "000000010",
                            2915 => "101110110",
                            2916 => "011101110",
                            2917 => "001011010",
                            2918 => "101000110",
                            2919 => "110001100",
                            2920 => "000011110",
                            2921 => "001010110",
                            2922 => "100011010",
                            2923 => "110011000",
                            2924 => "010100000",
                            2925 => "000100000",
                            2926 => "000000100",
                            2927 => "000000000",
                            2928 => "111000010",
                            2929 => "010011110",
                            2930 => "000000000",
                            2931 => "000000000",
                            2932 => "100111000",
                            2933 => "101101100",
                            2934 => "110100000",
                            2935 => "000101110",
                            2936 => "010010110",
                            2937 => "000010010",
                            2938 => "000000000",
                            2939 => "001001110",
                            2940 => "100100000",
                            2941 => "111001100",
                            2942 => "001000010",
                            2943 => "010101110",
                            2944 => "000010000",
                            2945 => "000000000",
                            2946 => "010001011",
                            2947 => "000000000",
                            2948 => "000000110",
                            2949 => "010100110",
                            2950 => "110111000",
                            2951 => "010011110",
                            2952 => "010000000",
                            2953 => "000000000",
                            2954 => "001101000",
                            2955 => "000001100",
                            2956 => "001110110",
                            2957 => "100011110",
                            2958 => "101000100",
                            2959 => "100111110",
                            2960 => "100010000",
                            2961 => "111010100",
                            2962 => "000010100",
                            2963 => "110100010",
                            2964 => "111101010",
                            2965 => "011010110",
                            2966 => "000000010",
                            2967 => "101110110",
                            2968 => "111001110",
                            2969 => "000101110",
                            2970 => "000011110",
                            2971 => "001010110",
                            2972 => "100011010",
                            2973 => "110011000",
                            2974 => "011101110",
                            2975 => "001011010",
                            2976 => "101000110",
                            2977 => "110001100",
                            2978 => "010100000",
                            2979 => "000110000",
                            2980 => "000000000",
                            2981 => "010101000",
                            2982 => "010000010",
                            2983 => "011011010",
                            2984 => "000000000",
                            2985 => "000000000",
                            2986 => "000101110",
                            2987 => "000000110",
                            2988 => "000000110",
                            2989 => "000000110",
                            2990 => "001001100",
                            2991 => "010010100",
                            2992 => "110111100",
                            2993 => "011011000",
                            2994 => "111000110",
                            2995 => "100110010",
                            2996 => "010111000",
                            2997 => "100001000",
                            2998 => "000111000",
                            2999 => "001011000",
                            3000 => "011011100",
                            3001 => "100011110",
                            3002 => "110100110",
                            3003 => "101101110",
                            3004 => "011111010",
                            3005 => "101111110",
                            3006 => "010000010",
                            3007 => "001101010",
                            3008 => "011001100",
                            3009 => "101111100",
                            3010 => "100001110",
                            3011 => "110001110",
                            3012 => "010111010",
                            3013 => "010111100",
                            3014 => "100010100",
                            3015 => "101010100",
                            3016 => "010010100",
                            3017 => "100010010",
                            3018 => "011000110",
                            3019 => "110111000",
                            3020 => "000100010",
                            3021 => "111010110",
                            3022 => "100010000",
                            3023 => "111110000",
                            3024 => "110100010",
                            3025 => "010011110",
                            3026 => "101111010",
                            3027 => "001111000",
                            3028 => "010111100",
                            3029 => "100101110",
                            3030 => "111100100",
                            3031 => "001110110",
                            3032 => "100111010",
                            3033 => "000001010",
                            3034 => "101000000",
                            3035 => "011111010",
                            3036 => "000110000",
                            3037 => "100001100",
                            3038 => "000011110",
                            3039 => "101010000",
                            3040 => "110100000",
                            3041 => "001000110",
                            3042 => "100111000",
                            3043 => "010110000",
                            3044 => "001010100",
                            3045 => "001011110",
                            3046 => "010100110",
                            3047 => "001101010",
                            3048 => "100101000",
                            3049 => "111100100",
                            3050 => "011011100",
                            3051 => "000010110",
                            3052 => "110101100",
                            3053 => "100100000",
                            3054 => "001011010",
                            3055 => "000111000",
                            3056 => "110111110",
                            3057 => "101100100",
                            3058 => "001100000",
                            3059 => "100101000",
                            3060 => "100010010",
                            3061 => "001010110",
                            3062 => "011010010",
                            3063 => "000110000",
                            3064 => "111110010",
                            3065 => "111111100",
                            3066 => "001000100",
                            3067 => "100110100",
                            3068 => "111000000",
                            3069 => "001101000",
                            3070 => "110111000",
                            3071 => "111010110",
                            3072 => "010110100",
                            3073 => "010100110",
                            3074 => "101010010",
                            3075 => "110000110",
                            3076 => "011110000",
                            3077 => "101101110",
                            3078 => "101001110",
                            3079 => "110000110",
                            3080 => "001110110",
                            3081 => "001110010",
                            3082 => "001111100",
                            3083 => "000100000",
                            3084 => "001101000",
                            3085 => "111000110",
                            3086 => "000000000",
                            3087 => "111010110",
                            3088 => "100011100",
                            3089 => "000000010",
                            3090 => "001011000",
                            3091 => "101001110",
                            3092 => "100010010",
                            3093 => "110100110",
                            3094 => "001000100",
                            3095 => "000011000",
                            3096 => "000111100",
                            3097 => "101101110",
                            3098 => "111000000",
                            3099 => "011100110",
                            3100 => "011000100",
                            3101 => "111100000",
                            3102 => "010001100",
                            3103 => "000001010",
                            3104 => "011001010",
                            3105 => "001001000",
                            3106 => "101111110",
                            3107 => "100000110",
                            3108 => "110010110",
                            3109 => "010110110",
                            3110 => "110000110",
                            3111 => "000010010",
                            3112 => "100101110",
                            3113 => "001011000",
                            3114 => "010100000",
                            3115 => "111110000",
                            3116 => "100001010",
                            3117 => "101010110",
                            3118 => "110101000",
                            3119 => "111001010",
                            3120 => "101000000",
                            3121 => "001011000",
                            3122 => "000010010",
                            3123 => "111110100",
                            3124 => "111011010",
                            3125 => "010011000",
                            3126 => "101100110",
                            3127 => "110111110",
                            3128 => "000101010",
                            3129 => "100111100",
                            3130 => "011011010",
                            3131 => "010100110",
                            3132 => "000110110",
                            3133 => "100011000",
                            3134 => "011100110",
                            3135 => "010000010",
                            3136 => "000010110",
                            3137 => "011000010",
                            3138 => "010110000",
                            3139 => "100110100",
                            3140 => "101011110",
                            3141 => "010111100",
                            3142 => "101100110",
                            3143 => "000010100",
                            3144 => "000000100",
                            3145 => "110101010",
                            3146 => "101000010",
                            3147 => "001000000",
                            3148 => "010110000",
                            3149 => "000001110",
                            3150 => "100000000",
                            3151 => "000111010",
                            3152 => "011110100",
                            3153 => "111000110",
                            3154 => "011111100",
                            3155 => "001000010",
                            3156 => "000100000",
                            3157 => "100001110",
                            3158 => "000101000",
                            3159 => "110000010",
                            3160 => "101011010",
                            3161 => "001010100",
                            3162 => "101111100",
                            3163 => "111111010",
                            3164 => "110111110",
                            3165 => "001111010",
                            3166 => "010001010",
                            3167 => "000010000",
                            3168 => "111011010",
                            3169 => "001110110",
                            3170 => "100111010",
                            3171 => "011001110",
                            3172 => "110110000",
                            3173 => "111110010",
                            3174 => "010110010",
                            3175 => "100110010",
                            3176 => "001001100",
                            3177 => "001111100",
                            3178 => "111001010",
                            3179 => "010110100",
                            3180 => "000000010",
                            3181 => "010111000",
                            3182 => "111100110",
                            3183 => "001111000",
                            3184 => "110101010",
                            3185 => "101011110",
                            3186 => "011110000",
                            3187 => "010100100",
                            3188 => "100001100",
                            3189 => "010101010",
                            3190 => "111101100",
                            3191 => "011011110",
                            3192 => "000011010",
                            3193 => "110100100",
                            3194 => "010101010",
                            3195 => "100011000",
                            3196 => "111011110",
                            3197 => "001110010",
                            3198 => "100100010",
                            3199 => "000001000",
                            3200 => "111000010",
                            3201 => "000010000",
                            3202 => "001010000",
                            3203 => "010101100",
                            3204 => "100001110",
                            3205 => "011100110",
                            3206 => "000010110",
                            3207 => "110110000",
                            3208 => "000101010",
                            3209 => "111000010",
                            3210 => "110001010",
                            3211 => "111110100",
                            3212 => "011110110",
                            3213 => "111001110",
                            3214 => "111011000",
                            3215 => "100000110",
                            3216 => "010010010",
                            3217 => "111111100",
                            3218 => "101010000",
                            3219 => "001010000",
                            3220 => "001100000",
                            3221 => "011100010",
                            3222 => "100011000",
                            3223 => "111111110",
                            3224 => "111011010",
                            3225 => "111111100",
                            3226 => "001001100",
                            3227 => "011000000",
                            3228 => "010100000",
                            3229 => "001100110",
                            3230 => "001000110",
                            3231 => "011101010",
                            3232 => "001010010",
                            3233 => "010110010",
                            3234 => "000110000",
                            3235 => "100111010",
                            3236 => "010111100",
                            3237 => "000010110",
                            3238 => "001000000",
                            3239 => "001000010",
                            3240 => "100111100",
                            3241 => "000111110",
                            3242 => "000011100",
                            3243 => "000100110",
                            3244 => "011010010",
                            3245 => "111111110",
                            3246 => "111011010",
                            3247 => "111100100",
                            3248 => "011001000",
                            3249 => "011000100",
                            3250 => "101111010",
                            3251 => "111111110",
                            3252 => "111100100",
                            3253 => "101010000",
                            3254 => "110001010",
                            3255 => "111011000",
                            3256 => "100110010",
                            3257 => "000001100",
                            3258 => "110111010",
                            3259 => "010011000",
                            3260 => "111011110",
                            3261 => "001100010",
                            3262 => "000011010",
                            3263 => "000100100",
                            3264 => "100011000",
                            3265 => "111010000",
                            3266 => "000110010",
                            3267 => "110101010",
                            3268 => "000100110",
                            3269 => "110100000",
                            3270 => "010110110",
                            3271 => "001010000",
                            3272 => "000110000",
                            3273 => "110101110",
                            3274 => "010111000",
                            3275 => "011111110",
                            3276 => "011010100",
                            3277 => "101001000",
                            3278 => "001110010",
                            3279 => "000110000",
                            3280 => "000101010",
                            3281 => "010010100",
                            3282 => "011010110",
                            3283 => "010010110",
                            3284 => "011101100",
                            3285 => "101000100",
                            3286 => "000110000",
                            3287 => "110001100",
                            3288 => "001100110",
                            3289 => "101101000",
                            3290 => "000010100",
                            3291 => "000010110",
                            3292 => "111011000",
                            3293 => "100010000",
                            3294 => "000111100",
                            3295 => "110111010",
                            3296 => "101111010",
                            3297 => "010001000",
                            3298 => "000111010",
                            3299 => "101010100",
                            3300 => "110011010",
                            3301 => "011001010",
                            3302 => "011001000",
                            3303 => "000101110",
                            3304 => "001001100",
                            3305 => "011001000",
                            3306 => "110100000",
                            3307 => "110000000",
                            3308 => "100110110",
                            3309 => "101100010",
                            3310 => "100011110",
                            3311 => "100101110",
                            3312 => "011000000",
                            3313 => "001010000",
                            3314 => "001000000",
                            3315 => "101100010",
                            3316 => "001011010",
                            3317 => "001011100",
                            3318 => "110011110",
                            3319 => "010010000",
                            3320 => "101000010",
                            3321 => "000011100",
                            3322 => "100100010",
                            3323 => "110110110",
                            3324 => "111001010",
                            3325 => "110111010",
                            3326 => "000111000",
                            3327 => "110101010",
                            3328 => "111011100",
                            3329 => "010100000",
                            3330 => "101101110",
                            3331 => "011010110",
                            3332 => "011010000",
                            3333 => "011110000",
                            3334 => "111110110",
                            3335 => "111100100",
                            3336 => "101010000",
                            3337 => "011010110",
                            3338 => "001101010",
                            3339 => "010110000",
                            3340 => "111010110",
                            3341 => "101101000",
                            3342 => "111101010",
                            3343 => "111101100",
                            3344 => "110100000",
                            3345 => "011001000",
                            3346 => "011110110",
                            3347 => "100010110",
                            3348 => "110001000",
                            3349 => "011010110",
                            3350 => "000100110",
                            3351 => "101001000",
                            3352 => "110110100",
                            3353 => "100111110",
                            3354 => "100101000",
                            3355 => "100010110",
                            3356 => "101100100",
                            3357 => "000101110",
                            3358 => "101111010",
                            3359 => "001111000",
                            3360 => "100000000",
                            3361 => "011100100",
                            3362 => "110111100",
                            3363 => "100110010",
                            3364 => "111000010",
                            3365 => "110101110",
                            3366 => "000010010",
                            3367 => "000010100",
                            3368 => "111100110",
                            3369 => "101001110",
                            3370 => "101110000",
                            3371 => "111010100",
                            3372 => "000011110",
                            3373 => "100000010",
                            3374 => "001101000",
                            3375 => "000101110",
                            3376 => "100010110",
                            3377 => "011001010",
                            3378 => "111001000",
                            3379 => "010011100",
                            3380 => "111111100",
                            3381 => "110101010",
                            3382 => "111001010",
                            3383 => "001100010",
                            3384 => "100000110",
                            3385 => "001110000",
                            3386 => "001111110",
                            3387 => "101111110",
                            3388 => "011100010",
                            3389 => "011110000",
                            3390 => "100001010",
                            3391 => "010011100",
                            3392 => "111101100",
                            3393 => "100111100",
                            3394 => "101010010",
                            3395 => "110111010",
                            3396 => "000110110",
                            3397 => "011010010",
                            3398 => "010011110",
                            3399 => "010010110",
                            3400 => "101011000",
                            3401 => "100010010",
                            3402 => "000111110",
                            3403 => "111001100",
                            3404 => "000011110",
                            3405 => "000011000",
                            3406 => "100000000",
                            3407 => "000100010",
                            3408 => "100001000",
                            3409 => "000111100",
                            3410 => "111001100",
                            3411 => "101011000",
                            3412 => "110101010",
                            3413 => "001111010",
                            3414 => "101111010",
                            3415 => "100110000",
                            3416 => "001111100",
                            3417 => "010001010",
                            3418 => "000110010",
                            3419 => "100011010",
                            3420 => "000101010",
                            3421 => "111010010",
                            3422 => "001101110",
                            3423 => "001011010",
                            3424 => "000101010",
                            3425 => "110000000",
                            3426 => "101100110",
                            3427 => "010000100",
                            3428 => "001110000",
                            3429 => "001000110",
                            3430 => "010110110",
                            3431 => "001011010",
                            3432 => "000011100",
                            3433 => "011110100",
                            3434 => "000100110",
                            3435 => "010111010",
                            3436 => "110011010",
                            3437 => "111011000",
                            3438 => "111011000",
                            3439 => "110011110",
                            3440 => "100110100",
                            3441 => "000100110",
                            3442 => "101101100",
                            3443 => "010000110",
                            3444 => "100111000",
                            3445 => "111111000",
                            3446 => "011001100",
                            3447 => "111000000",
                            3448 => "101011000",
                            3449 => "011010100",
                            3450 => "111101100",
                            3451 => "010100100",
                            3452 => "000100010",
                            3453 => "101100110",
                            3454 => "001010100",
                            3455 => "001011010",
                            3456 => "010110010",
                            3457 => "101100000",
                            3458 => "010000110",
                            3459 => "110010010",
                            3460 => "010101010",
                            3461 => "111011110",
                            3462 => "111001100",
                            3463 => "000001110",
                            3464 => "000001110",
                            3465 => "110101100",
                            3466 => "001010100",
                            3467 => "011101110",
                            3468 => "101101110",
                            3469 => "000001010",
                            3470 => "000000010",
                            3471 => "010101100",
                            3472 => "110100100",
                            3473 => "100110100",
                            3474 => "010000000",
                            3475 => "011000110",
                            3476 => "111000100",
                            3477 => "100100110",
                            3478 => "101000110",
                            3479 => "101000000",
                            3480 => "001000110",
                            3481 => "101110110",
                            3482 => "101001010",
                            3483 => "001100110",
                            3484 => "101001100",
                            3485 => "010101110",
                            3486 => "110001110",
                            3487 => "010111010",
                            3488 => "011001100",
                            3489 => "111111110",
                            3490 => "110110000",
                            3491 => "110111010",
                            3492 => "110110100",
                            3493 => "111100010",
                            3494 => "100111010",
                            3495 => "111110100",
                            3496 => "001011010",
                            3497 => "001110000",
                            3498 => "010100100",
                            3499 => "100101000",
                            3500 => "010110110",
                            3501 => "010110010",
                            3502 => "111110000",
                            3503 => "011110010",
                            3504 => "010010100",
                            3505 => "111101100",
                            3506 => "011010010",
                            3507 => "110010100",
                            3508 => "010101000",
                            3509 => "100010110",
                            3510 => "101111010",
                            3511 => "001110010",
                            3512 => "100110000",
                            3513 => "101010000",
                            3514 => "000100010",
                            3515 => "101101010",
                            3516 => "011010000",
                            3517 => "101111000",
                            3518 => "010101110",
                            3519 => "111001010",
                            3520 => "110110100",
                            3521 => "000111010",
                            3522 => "011100000",
                            3523 => "100101110",
                            3524 => "101010010",
                            3525 => "111101110",
                            3526 => "101010100",
                            3527 => "111011100",
                            3528 => "100101000",
                            3529 => "110001010",
                            3530 => "001111010",
                            3531 => "111110010",
                            3532 => "111011010",
                            3533 => "000100110",
                            3534 => "111110110",
                            3535 => "000110000",
                            3536 => "000011100",
                            3537 => "011110000",
                            3538 => "110110000",
                            3539 => "110010100",
                            3540 => "100011000",
                            3541 => "101100110",
                            3542 => "010111000",
                            3543 => "001000010",
                            3544 => "100011110",
                            3545 => "000011100",
                            3546 => "011010000",
                            3547 => "111101110",
                            3548 => "100001110",
                            3549 => "101000000",
                            3550 => "110000000",
                            3551 => "000010100",
                            3552 => "010100000",
                            3553 => "100000100",
                            3554 => "011000100",
                            3555 => "110011100",
                            3556 => "011011010",
                            3557 => "110000110",
                            3558 => "011110000",
                            3559 => "111100110",
                            3560 => "011000100",
                            3561 => "111101010",
                            3562 => "110010010",
                            3563 => "000011100",
                            3564 => "011111010",
                            3565 => "100011000",
                            3566 => "101111000",
                            3567 => "110111010",
                            3568 => "101001100",
                            3569 => "100001100",
                            3570 => "111000110",
                            3571 => "010010110",
                            3572 => "100010010",
                            3573 => "001011000",
                            3574 => "100110100",
                            3575 => "001101000",
                            3576 => "000011110",
                            3577 => "000000000",
                            3578 => "000011100",
                            3579 => "111100010",
                            3580 => "110101100",
                            3581 => "011011000",
                            3582 => "111101110",
                            3583 => "101001100",
                            3584 => "111000100",
                            3585 => "011100010",
                            3586 => "010000110",
                            3587 => "101101100",
                            3588 => "011110100",
                            3589 => "010011010",
                            3590 => "000001000",
                            3591 => "011110100",
                            3592 => "011110010",
                            3593 => "011110000",
                            3594 => "110111100",
                            3595 => "100001100",
                            3596 => "110001110",
                            3597 => "110101100",
                            3598 => "100000110",
                            3599 => "100101110",
                            3600 => "110000010",
                            3601 => "011000100",
                            3602 => "100010100",
                            3603 => "110111100",
                            3604 => "010010110",
                            3605 => "000110000",
                            3606 => "110011110",
                            3607 => "001000010",
                            3608 => "011101100",
                            3609 => "111101010",
                            3610 => "001000000",
                            3611 => "010010100",
                            3612 => "001010010",
                            3613 => "110001100",
                            3614 => "001101100",
                            3615 => "110011100",
                            3616 => "110110100",
                            3617 => "010110110",
                            3618 => "101010110",
                            3619 => "010101100",
                            3620 => "011110010",
                            3621 => "100101000",
                            3622 => "001100110",
                            3623 => "011001100",
                            3624 => "010010010",
                            3625 => "100101110",
                            3626 => "101011010",
                            3627 => "011100100",
                            3628 => "001000100",
                            3629 => "101000000",
                            3630 => "111111010",
                            3631 => "111001000",
                            3632 => "011111110",
                            3633 => "011101100",
                            3634 => "110000000",
                            3635 => "101101100",
                            3636 => "001000100",
                            3637 => "010100110",
                            3638 => "111100110",
                            3639 => "010101110",
                            3640 => "011010000",
                            3641 => "110111010",
                            3642 => "000011000",
                            3643 => "010110110",
                            3644 => "101111100",
                            3645 => "010110100",
                            3646 => "011101010",
                            3647 => "010001010",
                            3648 => "000001110",
                            3649 => "001010110",
                            3650 => "100001010",
                            3651 => "000111000",
                            3652 => "010110110",
                            3653 => "011010010",
                            3654 => "001011100",
                            3655 => "010111000",
                            3656 => "011110000",
                            3657 => "000011100",
                            3658 => "000010110",
                            3659 => "100010100",
                            3660 => "000010110",
                            3661 => "101111000",
                            3662 => "001000100",
                            3663 => "111000010",
                            3664 => "010000100",
                            3665 => "001101110",
                            3666 => "001000100",
                            3667 => "101101010",
                            3668 => "001000110",
                            3669 => "000010110",
                            3670 => "001000000",
                            3671 => "000100100",
                            3672 => "011001110",
                            3673 => "111000000",
                            3674 => "101011110",
                            3675 => "001100100",
                            3676 => "110000010",
                            3677 => "111101000",
                            3678 => "110111010",
                            3679 => "100101000",
                            3680 => "101011100",
                            3681 => "110011000",
                            3682 => "100100000",
                            3683 => "101010100",
                            3684 => "011001100",
                            3685 => "101100010",
                            3686 => "110100100",
                            3687 => "110011100",
                            3688 => "101110010",
                            3689 => "000111110",
                            3690 => "001101000",
                            3691 => "001011100",
                            3692 => "110101000",
                            3693 => "001110010",
                            3694 => "111001010",
                            3695 => "001101010",
                            3696 => "100011010",
                            3697 => "001101100",
                            3698 => "001000100",
                            3699 => "010001010",
                            3700 => "100010100",
                            3701 => "111001010",
                            3702 => "100000010",
                            3703 => "101101010",
                            3704 => "001010010",
                            3705 => "001111010",
                            3706 => "000010110",
                            3707 => "111011000",
                            3708 => "100001100",
                            3709 => "101100000",
                            3710 => "100101000",
                            3711 => "001001100",
                            3712 => "011001000",
                            3713 => "011101110",
                            3714 => "111111100",
                            3715 => "010111100",
                            3716 => "111101110",
                            3717 => "100011100",
                            3718 => "010101110",
                            3719 => "100111110",
                            3720 => "011111110",
                            3721 => "001010000",
                            3722 => "001010010",
                            3723 => "010110110",
                            3724 => "011111000",
                            3725 => "010011110",
                            3726 => "111001100",
                            3727 => "011101000",
                            3728 => "010001010",
                            3729 => "000000010",
                            3730 => "000001010",
                            3731 => "111001010",
                            3732 => "010111000",
                            3733 => "110111010",
                            3734 => "000010100",
                            3735 => "110100010",
                            3736 => "100111000",
                            3737 => "111011010",
                            3738 => "101001100",
                            3739 => "100110010",
                            3740 => "011101010",
                            3741 => "101011110",
                            3742 => "011111100",
                            3743 => "010000000",
                            3744 => "010000110",
                            3745 => "101101110",
                            3746 => "101110000",
                            3747 => "010100110",
                            3748 => "111010010",
                            3749 => "000010100",
                            3750 => "010010100",
                            3751 => "111001110",
                            3752 => "100100100",
                            3753 => "111011010",
                            3754 => "101011110",
                            3755 => "110000000",
                            3756 => "100110110",
                            3757 => "110000010",
                            3758 => "111101000",
                            3759 => "001011110",
                            3760 => "101011000",
                            3761 => "110000110",
                            3762 => "001111110",
                            3763 => "000011010",
                            3764 => "100010100",
                            3765 => "110010100",
                            3766 => "000000110",
                            3767 => "100101110",
                            3768 => "010011110",
                            3769 => "110010110",
                            3770 => "111000000",
                            3771 => "000001100",
                            3772 => "110011110",
                            3773 => "100100000",
                            3774 => "110010010",
                            3775 => "110111110",
                            3776 => "100101000",
                            3777 => "100001110",
                            3778 => "010100000",
                            3779 => "111000100",
                            3780 => "001010000",
                            3781 => "100010010",
                            3782 => "100001010",
                            3783 => "011110100",
                            3784 => "000111010",
                            3785 => "100101000",
                            3786 => "100001010",
                            3787 => "010110000",
                            3788 => "101001110",
                            3789 => "110111010",
                            3790 => "001100010",
                            3791 => "100101110",
                            3792 => "011000100",
                            3793 => "011001100",
                            3794 => "010111010",
                            3795 => "100100100",
                            3796 => "111011000",
                            3797 => "000000000",
                            3798 => "000000000",
                            3799 => "000011000",
                            3800 => "100111110",
                            3801 => "111100100",
                            3802 => "010101110",
                            3803 => "100111000",
                            3804 => "101101100",
                            3805 => "110100000",
                            3806 => "000101110",
                            3807 => "010010110",
                            3808 => "000010010",
                            3809 => "000010000",
                            3810 => "000000000",
                            3811 => "010001011",
                            3812 => "000000000",
                            3813 => "000000000",
                            3814 => "001010000",
                            3815 => "100101010",
                            3816 => "001100100",
                            3817 => "010000000",
                            3818 => "000000000",
                            3819 => "100000000",
                            3820 => "000001100",
                            3821 => "001110010",
                            3822 => "110101110",
                            3823 => "000010100",
                            3824 => "110100010",
                            3825 => "111101010",
                            3826 => "011010110",
                            3827 => "101000100",
                            3828 => "100111110",
                            3829 => "100010000",
                            3830 => "111010100",
                            3831 => "111001110",
                            3832 => "000101110",
                            3833 => "000000010",
                            3834 => "101110110",
                            3835 => "011101110",
                            3836 => "001011010",
                            3837 => "101000110",
                            3838 => "110001100",
                            3839 => "000011110",
                            3840 => "001010110",
                            3841 => "100100000",
                            3842 => "111101110",
                            3843 => "010100000",
                            3844 => "000100000",
                            3845 => "000000010",
                            3846 => "111111010",
                            3847 => "110111100",
                            3848 => "001001110",
                            3849 => "000000000",
                            3850 => "000000000",
                            3851 => "100111000",
                            3852 => "101101100",
                            3853 => "110100000",
                            3854 => "000101110",
                            3855 => "010010110",
                            3856 => "000010010",
                            3857 => "000000000",
                            3858 => "001001110",
                            3859 => "100100000",
                            3860 => "111001100",
                            3861 => "001000010",
                            3862 => "010101110",
                            3863 => "000010000",
                            3864 => "000000000",
                            3865 => "010001011",
                            3866 => "000000000",
                            3867 => "000000010",
                            3868 => "011001110",
                            3869 => "110111000",
                            3870 => "010100000",
                            3871 => "010000000",
                            3872 => "000000000",
                            3873 => "001101000",
                            3874 => "000001100",
                            3875 => "001111010",
                            3876 => "011110100",
                            3877 => "101000100",
                            3878 => "100111110",
                            3879 => "100010000",
                            3880 => "111010100",
                            3881 => "000010100",
                            3882 => "110100010",
                            3883 => "111101010",
                            3884 => "011010110",
                            3885 => "000000010",
                            3886 => "101110110",
                            3887 => "111001110",
                            3888 => "000101110",
                            3889 => "000011110",
                            3890 => "001010110",
                            3891 => "100100000",
                            3892 => "111101110",
                            3893 => "011101110",
                            3894 => "001011010",
                            3895 => "101000110",
                            3896 => "110001100",
                            3897 => "010100000",
                            3898 => "000110000",
                            3899 => "000000000",
                            3900 => "010101000",
                            3901 => "101001100",
                            3902 => "001010100",
                            3903 => "000000000",
                            3904 => "000000000",
                            3905 => "000101110",
                            3906 => "000000110",
                            3907 => "000000110",
                            3908 => "000000010",
                            3909 => "001110100",
                            3910 => "111110100",
                            3911 => "011101100",
                            3912 => "011100000",
                            3913 => "101111000",
                            3914 => "000101010",
                            3915 => "100011010",
                            3916 => "101010010",
                            3917 => "011011010",
                            3918 => "011111010",
                            3919 => "010000100",
                            3920 => "010000000",
                            3921 => "101101010",
                            3922 => "100110010",
                            3923 => "011001100",
                            3924 => "000011100",
                            3925 => "000001010",
                            3926 => "010010000",
                            3927 => "101000100",
                            3928 => "000000000",
                            3929 => "111010100",
                            3930 => "000110010",
                            3931 => "010000010",
                            3932 => "011110110",
                            3933 => "010011100",
                            3934 => "010110000",
                            3935 => "000100000",
                            3936 => "010001110",
                            3937 => "101000000",
                            3938 => "110111110",
                            3939 => "110111010",
                            3940 => "011111010",
                            3941 => "111000010",
                            3942 => "011111110",
                            3943 => "100111000",
                            3944 => "001100010",
                            3945 => "000110000",
                            3946 => "100011000",
                            3947 => "100011100",
                            3948 => "110011100",
                            3949 => "000100010",
                            3950 => "000111010",
                            3951 => "011001000",
                            3952 => "010011110",
                            3953 => "100110010",
                            3954 => "100101000",
                            3955 => "000000000",
                            3956 => "000101000",
                            3957 => "111100000",
                            3958 => "111000100",
                            3959 => "101101000",
                            3960 => "001111110",
                            3961 => "100000010",
                            3962 => "101000000",
                            3963 => "111001010",
                            3964 => "011100000",
                            3965 => "000011010",
                            3966 => "101001000",
                            3967 => "011100010",
                            3968 => "001101110",
                            3969 => "011010110",
                            3970 => "000110100",
                            3971 => "001100100",
                            3972 => "111101000",
                            3973 => "010011110",
                            3974 => "100111000",
                            3975 => "001001110",
                            3976 => "011010110",
                            3977 => "100000100",
                            3978 => "001101000",
                            3979 => "110010100",
                            3980 => "010100110",
                            3981 => "010101000",
                            3982 => "011111000",
                            3983 => "011000010",
                            3984 => "100011110",
                            3985 => "110110010",
                            3986 => "000011010",
                            3987 => "010001100",
                            3988 => "001111110",
                            3989 => "000101000",
                            3990 => "001001000",
                            3991 => "011001100",
                            3992 => "101000010",
                            3993 => "010101100",
                            3994 => "001010000",
                            3995 => "111110000",
                            3996 => "011111110",
                            3997 => "101100110",
                            3998 => "111000010",
                            3999 => "100010110",
                            4000 => "111111000",
                            4001 => "000100110",
                            4002 => "110001110",
                            4003 => "101101100",
                            4004 => "100111000",
                            4005 => "010101110",
                            4006 => "100101000",
                            4007 => "110000000",
                            4008 => "010001100",
                            4009 => "110100100",
                            4010 => "100100110",
                            4011 => "110111100",
                            4012 => "111110000",
                            4013 => "100001110",
                            4014 => "111110100",
                            4015 => "110100000",
                            4016 => "001100100",
                            4017 => "011100110",
                            4018 => "110001010",
                            4019 => "011101010",
                            4020 => "110111010",
                            4021 => "101010010",
                            4022 => "111100010",
                            4023 => "111110110",
                            4024 => "011101000",
                            4025 => "000111110",
                            4026 => "010010110",
                            4027 => "100100000",
                            4028 => "111100110",
                            4029 => "110010000",
                            4030 => "101011100",
                            4031 => "011110100",
                            4032 => "001100110",
                            4033 => "010110010",
                            4034 => "010100010",
                            4035 => "110011000",
                            4036 => "011100100",
                            4037 => "011110100",
                            4038 => "010111110",
                            4039 => "110110100",
                            4040 => "110101000",
                            4041 => "011010110",
                            4042 => "110010110",
                            4043 => "111101100",
                            4044 => "001010110",
                            4045 => "000110010",
                            4046 => "101101000",
                            4047 => "101101110",
                            4048 => "000100010",
                            4049 => "011111000",
                            4050 => "011010000",
                            4051 => "001110000",
                            4052 => "101110110",
                            4053 => "101000010",
                            4054 => "010111100",
                            4055 => "100101100",
                            4056 => "010000000",
                            4057 => "101110110",
                            4058 => "001001110",
                            4059 => "110010000",
                            4060 => "010101000",
                            4061 => "110110110",
                            4062 => "100011010",
                            4063 => "011000000",
                            4064 => "101011010",
                            4065 => "111011100",
                            4066 => "111110010",
                            4067 => "011100010",
                            4068 => "101000000",
                            4069 => "110011000",
                            4070 => "110001100",
                            4071 => "111010010",
                            4072 => "000101000",
                            4073 => "011110000",
                            4074 => "101001000",
                            4075 => "000111100",
                            4076 => "100011000",
                            4077 => "111100110",
                            4078 => "111000000",
                            4079 => "101100000",
                            4080 => "101001000",
                            4081 => "010110000",
                            4082 => "110010010",
                            4083 => "011101100",
                            4084 => "111101000",
                            4085 => "100000000",
                            4086 => "000110000",
                            4087 => "110010000",
                            4088 => "001010100",
                            4089 => "000101000",
                            4090 => "000010100",
                            4091 => "001000000",
                            4092 => "111111100",
                            4093 => "101011110",
                            4094 => "101011100",
                            4095 => "000111110",
                            4096 => "100011000",
                            4097 => "110111100",
                            4098 => "111011110",
                            4099 => "011001100",
                            4100 => "100111100",
                            4101 => "111010010",
                            4102 => "011010110",
                            4103 => "000011000",
                            4104 => "010010100",
                            4105 => "101010010",
                            4106 => "000111000",
                            4107 => "010001000",
                            4108 => "010111010",
                            4109 => "101001000",
                            4110 => "011110010",
                            4111 => "100111110",
                            4112 => "010110000",
                            4113 => "000100110",
                            4114 => "011110110",
                            4115 => "011001110",
                            4116 => "101010110",
                            4117 => "011001110",
                            4118 => "010111010",
                            4119 => "111011100",
                            4120 => "110000100",
                            4121 => "100101100",
                            4122 => "001001000",
                            4123 => "110111010",
                            4124 => "111011000",
                            4125 => "100001000",
                            4126 => "101110010",
                            4127 => "001001000",
                            4128 => "001011110",
                            4129 => "000100110",
                            4130 => "110110100",
                            4131 => "101011110",
                            4132 => "101101000",
                            4133 => "110001110",
                            4134 => "110100100",
                            4135 => "110100100",
                            4136 => "110111110",
                            4137 => "101010110",
                            4138 => "110101100",
                            4139 => "111100110",
                            4140 => "100011010",
                            4141 => "001110000",
                            4142 => "011000100",
                            4143 => "000111000",
                            4144 => "001110100",
                            4145 => "100100010",
                            4146 => "100000100",
                            4147 => "111001010",
                            4148 => "101010110",
                            4149 => "011000100",
                            4150 => "100111110",
                            4151 => "010110010",
                            4152 => "100111000",
                            4153 => "000111100",
                            4154 => "001010100",
                            4155 => "101111000",
                            4156 => "001111110",
                            4157 => "001110110",
                            4158 => "010100000",
                            4159 => "001100010",
                            4160 => "100000000",
                            4161 => "000000100",
                            4162 => "111110110",
                            4163 => "101000100",
                            4164 => "010000110",
                            4165 => "010010100",
                            4166 => "001011000",
                            4167 => "100010010",
                            4168 => "001011100",
                            4169 => "100101010",
                            4170 => "100101100",
                            4171 => "011101100",
                            4172 => "111001110",
                            4173 => "100001100",
                            4174 => "011010100",
                            4175 => "110110110",
                            4176 => "110000010",
                            4177 => "101100100",
                            4178 => "100111000",
                            4179 => "110001000",
                            4180 => "011110110",
                            4181 => "000001000",
                            4182 => "010101000",
                            4183 => "011011100",
                            4184 => "001110100",
                            4185 => "110111000",
                            4186 => "001000110",
                            4187 => "010010010",
                            4188 => "111100000",
                            4189 => "100111110",
                            4190 => "011001000",
                            4191 => "100110110",
                            4192 => "011011010",
                            4193 => "100111110",
                            4194 => "001010100",
                            4195 => "001001100",
                            4196 => "111110000",
                            4197 => "010001000",
                            4198 => "011010110",
                            4199 => "101001010",
                            4200 => "101111110",
                            4201 => "111001110",
                            4202 => "101000100",
                            4203 => "010100110",
                            4204 => "101110100",
                            4205 => "110100000",
                            4206 => "001101000",
                            4207 => "011010000",
                            4208 => "111101110",
                            4209 => "010011010",
                            4210 => "001100000",
                            4211 => "100101010",
                            4212 => "101011010",
                            4213 => "001101010",
                            4214 => "000011000",
                            4215 => "011100000",
                            4216 => "111111100",
                            4217 => "000110110",
                            4218 => "110101000",
                            4219 => "000011010",
                            4220 => "110000110",
                            4221 => "100011000",
                            4222 => "110101110",
                            4223 => "101101000",
                            4224 => "000000000",
                            4225 => "000000000",
                            4226 => "000011000",
                            4227 => "100111110",
                            4228 => "111100100",
                            4229 => "010101110",
                            4230 => "100111000",
                            4231 => "101101100",
                            4232 => "110100000",
                            4233 => "000101110",
                            4234 => "010010110",
                            4235 => "000010010",
                            4236 => "000010000",
                            4237 => "000000000",
                            4238 => "010001011",
                            4239 => "000000000",
                            4240 => "000000000",
                            4241 => "001010000",
                            4242 => "100101010",
                            4243 => "001100110",
                            4244 => "010000000",
                            4245 => "000000000",
                            4246 => "100000000",
                            4247 => "000001100",
                            4248 => "001110010",
                            4249 => "110101100",
                            4250 => "000010100",
                            4251 => "110100010",
                            4252 => "111101010",
                            4253 => "011010110",
                            4254 => "101000100",
                            4255 => "100111110",
                            4256 => "100010000",
                            4257 => "111010100",
                            4258 => "111001110",
                            4259 => "000101110",
                            4260 => "000000010",
                            4261 => "101110110",
                            4262 => "011101110",
                            4263 => "001011010",
                            4264 => "101000110",
                            4265 => "110001100",
                            4266 => "000011110",
                            4267 => "001010110",
                            4268 => "100100100",
                            4269 => "001101100",
                            4270 => "010100000",
                            4271 => "000100000",
                            4272 => "000000010",
                            4273 => "111111000",
                            4274 => "110111000",
                            4275 => "111010010",
                            4276 => "000000000",
                            4277 => "000000000",
                            4278 => "100111000",
                            4279 => "101101100",
                            4280 => "110100000",
                            4281 => "000101110",
                            4282 => "010010110",
                            4283 => "000010010",
                            4284 => "000000000",
                            4285 => "001001110",
                            4286 => "100100000",
                            4287 => "111001100",
                            4288 => "001000010",
                            4289 => "010101110",
                            4290 => "000010000",
                            4291 => "000000000",
                            4292 => "010001011",
                            4293 => "000000000",
                            4294 => "000000010",
                            4295 => "010101100",
                            4296 => "110111000",
                            4297 => "010100010",
                            4298 => "010000000",
                            4299 => "000000000",
                            4300 => "001101000",
                            4301 => "000001100",
                            4302 => "001111010",
                            4303 => "100010100",
                            4304 => "101000100",
                            4305 => "100111110",
                            4306 => "100010000",
                            4307 => "111010100",
                            4308 => "000010100",
                            4309 => "110100010",
                            4310 => "111101010",
                            4311 => "011010110",
                            4312 => "000000010",
                            4313 => "101110110",
                            4314 => "111001110",
                            4315 => "000101110",
                            4316 => "000011110",
                            4317 => "001010110",
                            4318 => "100100100",
                            4319 => "001101100",
                            4320 => "011101110",
                            4321 => "001011010",
                            4322 => "101000110",
                            4323 => "110001100",
                            4324 => "010100000",
                            4325 => "000110000",
                            4326 => "000000000",
                            4327 => "010101000",
                            4328 => "110001110",
                            4329 => "001100110",
                            4330 => "000000000",
                            4331 => "000000000",
                            4332 => "000101110",
                            4333 => "000000110",
                            4334 => "000000110",
                            4335 => "000000010",
                            4336 => "001010010",
                            4337 => "010010010",
                            4338 => "100000100",
                            4339 => "100011000",
                            4340 => "010111010",
                            4341 => "000111010",
                            4342 => "001101110",
                            4343 => "011001110",
                            4344 => "101000110",
                            4345 => "110000110",
                            4346 => "111101000",
                            4347 => "110111110",
                            4348 => "000010100",
                            4349 => "110100100",
                            4350 => "010101000",
                            4351 => "000001100",
                            4352 => "101101000",
                            4353 => "000101000",
                            4354 => "001010010",
                            4355 => "000100110",
                            4356 => "110001110",
                            4357 => "111011000",
                            4358 => "001011010",
                            4359 => "101010010",
                            4360 => "011010000",
                            4361 => "000000100",
                            4362 => "111011100",
                            4363 => "000110110",
                            4364 => "110101110",
                            4365 => "011001000",
                            4366 => "000111000",
                            4367 => "101100100",
                            4368 => "010010110",
                            4369 => "110100100",
                            4370 => "000011000",
                            4371 => "101111000",
                            4372 => "001101010",
                            4373 => "010011110",
                            4374 => "101110110",
                            4375 => "100000100",
                            4376 => "110101110",
                            4377 => "000100000",
                            4378 => "011000110",
                            4379 => "101011110",
                            4380 => "110001000",
                            4381 => "011000100",
                            4382 => "111111100",
                            4383 => "101001010",
                            4384 => "001011110",
                            4385 => "001010100",
                            4386 => "100000010",
                            4387 => "000111100",
                            4388 => "111110100",
                            4389 => "010100010",
                            4390 => "111010110",
                            4391 => "000111010",
                            4392 => "100110000",
                            4393 => "011000100",
                            4394 => "111110110",
                            4395 => "101110110",
                            4396 => "001001000",
                            4397 => "011011000",
                            4398 => "011111000",
                            4399 => "000111000",
                            4400 => "011010000",
                            4401 => "000110100",
                            4402 => "111011010",
                            4403 => "100111100",
                            4404 => "001111000",
                            4405 => "111111110",
                            4406 => "100000010",
                            4407 => "110100100",
                            4408 => "001101000",
                            4409 => "000011110",
                            4410 => "101101110",
                            4411 => "011101100",
                            4412 => "000110110",
                            4413 => "010010100",
                            4414 => "100011000",
                            4415 => "110000010",
                            4416 => "100101110",
                            4417 => "100101000",
                            4418 => "100101100",
                            4419 => "001000010",
                            4420 => "110001000",
                            4421 => "011101100",
                            4422 => "010110010",
                            4423 => "011100000",
                            4424 => "111000000",
                            4425 => "101011010",
                            4426 => "101001100",
                            4427 => "001100110",
                            4428 => "000111100",
                            4429 => "001100110",
                            4430 => "010110110",
                            4431 => "001001010",
                            4432 => "010111100",
                            4433 => "011011100",
                            4434 => "101001100",
                            4435 => "110011000",
                            4436 => "000000010",
                            4437 => "110101100",
                            4438 => "100111000",
                            4439 => "100011100",
                            4440 => "111101010",
                            4441 => "000100000",
                            4442 => "111011100",
                            4443 => "100110010",
                            4444 => "011010100",
                            4445 => "010110110",
                            4446 => "010001110",
                            4447 => "111000110",
                            4448 => "010011100",
                            4449 => "100111110",
                            4450 => "111111010",
                            4451 => "000001000",
                            4452 => "010110000",
                            4453 => "011110010",
                            4454 => "100011000",
                            4455 => "011000010",
                            4456 => "001101000",
                            4457 => "000000110",
                            4458 => "000000100",
                            4459 => "010101010",
                            4460 => "000010010",
                            4461 => "011000110",
                            4462 => "111001010",
                            4463 => "010100110",
                            4464 => "111111000",
                            4465 => "001010100",
                            4466 => "010110110",
                            4467 => "110000000",
                            4468 => "111001100",
                            4469 => "011100010",
                            4470 => "001100110",
                            4471 => "010101110",
                            4472 => "001101110",
                            4473 => "000110110",
                            4474 => "011101110",
                            4475 => "010100000",
                            4476 => "111001100",
                            4477 => "000000110",
                            4478 => "010010100",
                            4479 => "110100000",
                            4480 => "100000100",
                            4481 => "000000000",
                            4482 => "011000010",
                            4483 => "000010100",
                            4484 => "110000010",
                            4485 => "111000000",
                            4486 => "001101110",
                            4487 => "001110100",
                            4488 => "100010100",
                            4489 => "000010000",
                            4490 => "011111110",
                            4491 => "011100000",
                            4492 => "001010010",
                            4493 => "000101000",
                            4494 => "111001100",
                            4495 => "100011000",
                            4496 => "111110000",
                            4497 => "010100010",
                            4498 => "010010000",
                            4499 => "010111100",
                            4500 => "100011100",
                            4501 => "101011110",
                            4502 => "110110010",
                            4503 => "110110100",
                            4504 => "110000110",
                            4505 => "110110010",
                            4506 => "110011010",
                            4507 => "110101000",
                            4508 => "011011100",
                            4509 => "100101110",
                            4510 => "101110010",
                            4511 => "111100110",
                            4512 => "111111010",
                            4513 => "111101010",
                            4514 => "111111000",
                            4515 => "111001100",
                            4516 => "101011110",
                            4517 => "001011110",
                            4518 => "011110000",
                            4519 => "100001010",
                            4520 => "110111000",
                            4521 => "101100100",
                            4522 => "111111000",
                            4523 => "101010010",
                            4524 => "110111000",
                            4525 => "010110010",
                            4526 => "001001110",
                            4527 => "111110110",
                            4528 => "001100010",
                            4529 => "101000100",
                            4530 => "000100110",
                            4531 => "111001010",
                            4532 => "110001000",
                            4533 => "001111100",
                            4534 => "111101000",
                            4535 => "100100100",
                            4536 => "111111110",
                            4537 => "100010000",
                            4538 => "101000110",
                            4539 => "000011100",
                            4540 => "100000000",
                            4541 => "000010110",
                            4542 => "010101110",
                            4543 => "110000000",
                            4544 => "111100010",
                            4545 => "011100000",
                            4546 => "101111000",
                            4547 => "111111100",
                            4548 => "001011010",
                            4549 => "111011100",
                            4550 => "101101100",
                            4551 => "110001010",
                            4552 => "010101110",
                            4553 => "110000010",
                            4554 => "110100110",
                            4555 => "110010010",
                            4556 => "000111000",
                            4557 => "101110010",
                            4558 => "100001110",
                            4559 => "110010000",
                            4560 => "000100010",
                            4561 => "000100000",
                            4562 => "000110010",
                            4563 => "100010000",
                            4564 => "011110000",
                            4565 => "011000100",
                            4566 => "011001110",
                            4567 => "000111010",
                            4568 => "000101100",
                            4569 => "001100010",
                            4570 => "111011100",
                            4571 => "001001000",
                            4572 => "111101110",
                            4573 => "011110000",
                            4574 => "110001000",
                            4575 => "111010010",
                            4576 => "000101100",
                            4577 => "101011010",
                            4578 => "011001000",
                            4579 => "010111110",
                            4580 => "100101000",
                            4581 => "001101100",
                            4582 => "100101110",
                            4583 => "000010010",
                            4584 => "001000010",
                            4585 => "100000110",
                            4586 => "001000000",
                            4587 => "111111010",
                            4588 => "110000010",
                            4589 => "010100000",
                            4590 => "101011010",
                            4591 => "111010000",
                            4592 => "001100010",
                            4593 => "111010010",
                            4594 => "110001010",
                            4595 => "110001010",
                            4596 => "110001000",
                            4597 => "000100000",
                            4598 => "011001100",
                            4599 => "101100010",
                            4600 => "101000000",
                            4601 => "100000100",
                            4602 => "000001110",
                            4603 => "010001100",
                            4604 => "000000100",
                            4605 => "011001100",
                            4606 => "110111010",
                            4607 => "000001000",
                            4608 => "001100010",
                            4609 => "010100010",
                            4610 => "111011000",
                            4611 => "010100000",
                            4612 => "010010110",
                            4613 => "001110010",
                            4614 => "010110010",
                            4615 => "001100000",
                            4616 => "001001010",
                            4617 => "000100010",
                            4618 => "010000100",
                            4619 => "101100000",
                            4620 => "011110010",
                            4621 => "001110110",
                            4622 => "000100010",
                            4623 => "000011010",
                            4624 => "010001100",
                            4625 => "110000110",
                            4626 => "101000110",
                            4627 => "110111000",
                            4628 => "111111100",
                            4629 => "000010010",
                            4630 => "000110110",
                            4631 => "101110000",
                            4632 => "000001110",
                            4633 => "111110010",
                            4634 => "000000000",
                            4635 => "000000000",
                            4636 => "000011000",
                            4637 => "100111110",
                            4638 => "111100100",
                            4639 => "010101110",
                            4640 => "100111000",
                            4641 => "101101100",
                            4642 => "110100000",
                            4643 => "000101110",
                            4644 => "010010110",
                            4645 => "000010010",
                            4646 => "000010000",
                            4647 => "000000000",
                            4648 => "010001011",
                            4649 => "000000000",
                            4650 => "000000000",
                            4651 => "001010000",
                            4652 => "100101010",
                            4653 => "001101000",
                            4654 => "010000000",
                            4655 => "000000000",
                            4656 => "100000000",
                            4657 => "000001100",
                            4658 => "001110010",
                            4659 => "110101010",
                            4660 => "000010100",
                            4661 => "110100010",
                            4662 => "111101010",
                            4663 => "011010110",
                            4664 => "101000100",
                            4665 => "100111110",
                            4666 => "100010000",
                            4667 => "111010100",
                            4668 => "111001110",
                            4669 => "000101110",
                            4670 => "000000010",
                            4671 => "101110110",
                            4672 => "011101110",
                            4673 => "001011010",
                            4674 => "101000110",
                            4675 => "110001100",
                            4676 => "000011110",
                            4677 => "001010110",
                            4678 => "100100110",
                            4679 => "011001000",
                            4680 => "010100000",
                            4681 => "000100000",
                            4682 => "000000100",
                            4683 => "000000000",
                            4684 => "110110110",
                            4685 => "101101110",
                            4686 => "000000000",
                            4687 => "000000000",
                            4688 => "100111000",
                            4689 => "101101100",
                            4690 => "110100000",
                            4691 => "000101110",
                            4692 => "010010110",
                            4693 => "000010010",
                            4694 => "000000000",
                            4695 => "001001110",
                            4696 => "100100000",
                            4697 => "111001100",
                            4698 => "001000010",
                            4699 => "010101110",
                            4700 => "000010000",
                            4701 => "000000000",
                            4702 => "010001011",
                            4703 => "000000000",
                            4704 => "000000000",
                            4705 => "011110110",
                            4706 => "110111000",
                            4707 => "010100100",
                            4708 => "010000000",
                            4709 => "000000000",
                            4710 => "001101000",
                            4711 => "000001100",
                            4712 => "001111100",
                            4713 => "011001000",
                            4714 => "101000100",
                            4715 => "100111110",
                            4716 => "100010000",
                            4717 => "111010100",
                            4718 => "000010100",
                            4719 => "110100010",
                            4720 => "111101010",
                            4721 => "011010110",
                            4722 => "000000010",
                            4723 => "101110110",
                            4724 => "111001110",
                            4725 => "000101110",
                            4726 => "000011110",
                            4727 => "001010110",
                            4728 => "100100110",
                            4729 => "011001000",
                            4730 => "011101110",
                            4731 => "001011010",
                            4732 => "101000110",
                            4733 => "110001100",
                            4734 => "010100000",
                            4735 => "000110000",
                            4736 => "000000000",
                            4737 => "010101000",
                            4738 => "001000110",
                            4739 => "111000010",
                            4740 => "000000000",
                            4741 => "000000000",
                            4742 => "000101110",
                            4743 => "000000110",
                            4744 => "000000110",
                            4745 => "000000000",
                            4746 => "010011100",
                            4747 => "010000100",
                            4748 => "001000100",
                            4749 => "000000100",
                            4750 => "000001010",
                            4751 => "110101000",
                            4752 => "101111110",
                            4753 => "000101110",
                            4754 => "010001110",
                            4755 => "001011010",
                            4756 => "011101000",
                            4757 => "110001000",
                            4758 => "100100110",
                            4759 => "100100110",
                            4760 => "110000110",
                            4761 => "100000010",
                            4762 => "011111100",
                            4763 => "100101100",
                            4764 => "001101000",
                            4765 => "101111110",
                            4766 => "001110000",
                            4767 => "100100010",
                            4768 => "110011010",
                            4769 => "011010000",
                            4770 => "110111110",
                            4771 => "000110100",
                            4772 => "110001010",
                            4773 => "010100000",
                            4774 => "101111100",
                            4775 => "011000100",
                            4776 => "101101000",
                            4777 => "100101110",
                            4778 => "111110110",
                            4779 => "110010100",
                            4780 => "101011100",
                            4781 => "000011100",
                            4782 => "101101110",
                            4783 => "111111000",
                            4784 => "001010100",
                            4785 => "001100110",
                            4786 => "110000000",
                            4787 => "001100110",
                            4788 => "100001010",
                            4789 => "000101100",
                            4790 => "011001000",
                            4791 => "111001010",
                            4792 => "110101010",
                            4793 => "111010100",
                            4794 => "100011000",
                            4795 => "011111100",
                            4796 => "111010010",
                            4797 => "101110000",
                            4798 => "101011110",
                            4799 => "000001010",
                            4800 => "000101110",
                            4801 => "011011110",
                            4802 => "011100000",
                            4803 => "001110000",
                            4804 => "001001010",
                            4805 => "000111110",
                            4806 => "100100010",
                            4807 => "110011100",
                            4808 => "100100100",
                            4809 => "001111010",
                            4810 => "000111100",
                            4811 => "110101000",
                            4812 => "001001000",
                            4813 => "110001000",
                            4814 => "101111110",
                            4815 => "000011000",
                            4816 => "111010100",
                            4817 => "000010100",
                            4818 => "010100000",
                            4819 => "111101100",
                            4820 => "111010000",
                            4821 => "000111010",
                            4822 => "100010100",
                            4823 => "001111100",
                            4824 => "110101000",
                            4825 => "000000000",
                            4826 => "000000000",
                            4827 => "000011000",
                            4828 => "100111110",
                            4829 => "111100100",
                            4830 => "010101110",
                            4831 => "100111000",
                            4832 => "101101100",
                            4833 => "110100000",
                            4834 => "000101110",
                            4835 => "010010110",
                            4836 => "000010010",
                            4837 => "000010000",
                            4838 => "000000000",
                            4839 => "010001011",
                            4840 => "000000000",
                            4841 => "000000000",
                            4842 => "001010000",
                            4843 => "100101010",
                            4844 => "001101010",
                            4845 => "010000000",
                            4846 => "000000000",
                            4847 => "100000000",
                            4848 => "000001100",
                            4849 => "001110010",
                            4850 => "110101000",
                            4851 => "000010100",
                            4852 => "110100010",
                            4853 => "111101010",
                            4854 => "011010110",
                            4855 => "101000100",
                            4856 => "100111110",
                            4857 => "100010000",
                            4858 => "111010100",
                            4859 => "111001110",
                            4860 => "000101110",
                            4861 => "000000010",
                            4862 => "101110110",
                            4863 => "011101110",
                            4864 => "001011010",
                            4865 => "101000110",
                            4866 => "110001100",
                            4867 => "000011110",
                            4868 => "001010110",
                            4869 => "100100110",
                            4870 => "101101110",
                            4871 => "010100000",
                            4872 => "000100000",
                            4873 => "000000100",
                            4874 => "000000000",
                            4875 => "110110110",
                            4876 => "011001000",
                            4877 => "000000000",
                            4878 => "000000000",
                            4879 => "100111000",
                            4880 => "101101100",
                            4881 => "110100000",
                            4882 => "000101110",
                            4883 => "010010110",
                            4884 => "000010010",
                            4885 => "000000000",
                            4886 => "001001110",
                            4887 => "100100000",
                            4888 => "111001100",
                            4889 => "001000010",
                            4890 => "010101110",
                            4891 => "000010000",
                            4892 => "000000000",
                            4893 => "010001011",
                            4894 => "000000000",
                            4895 => "000000010",
                            4896 => "111011110",
                            4897 => "111000000",
                            4898 => "011001010",
                            4899 => "000000000",
                            4900 => "000000000",
                            4901 => "001101000",
                            4902 => "000001100",
                            4903 => "110101100",
                            4904 => "001011010",
                            4905 => "010010100",
                            4906 => "011111010",
                            4907 => "100000110",
                            4908 => "101111000",
                            4909 => "000010100",
                            4910 => "110100010",
                            4911 => "111101010",
                            4912 => "011010110",
                            4913 => "000101000",
                            4914 => "011011000",
                            4915 => "111001100",
                            4916 => "101011010",
                            4917 => "011000010",
                            4918 => "010111110",
                            4919 => "011000110",
                            4920 => "110001000",
                            4921 => "110100010",
                            4922 => "010111100",
                            4923 => "111110100",
                            4924 => "010101110",
                            4925 => "010100000",
                            4926 => "000110000",
                            4927 => "000000010",
                            4928 => "000010010",
                            4929 => "000010100",
                            4930 => "010000100",
                            4931 => "000000000",
                            4932 => "000000000",
                            4933 => "000101110",
                            4934 => "000000110",
                            4935 => "000000110",
                            4936 => "000000010",
                            4937 => "110000100",
                            4938 => "000001010",
                            4939 => "010101000",
                            4940 => "000000000",
                            4941 => "000011010",
                            4942 => "001110000",
                            4943 => "011000000",
                            4944 => "001010100",
                            4945 => "101011000",
                            4946 => "100010000",
                            4947 => "001101110",
                            4948 => "110000110",
                            4949 => "100100000",
                            4950 => "100110000",
                            4951 => "101001100",
                            4952 => "001010000",
                            4953 => "100101110",
                            4954 => "011111110",
                            4955 => "011011000",
                            4956 => "111100100",
                            4957 => "110001110",
                            4958 => "101000110",
                            4959 => "001100000",
                            4960 => "101110100",
                            4961 => "111110110",
                            4962 => "111100110",
                            4963 => "010001100",
                            4964 => "010010000",
                            4965 => "111010010",
                            4966 => "000011010",
                            4967 => "000001110",
                            4968 => "000010100",
                            4969 => "111111010",
                            4970 => "010111000",
                            4971 => "000011010",
                            4972 => "011000000",
                            4973 => "100100100",
                            4974 => "000100000",
                            4975 => "001000000",
                            4976 => "001111110",
                            4977 => "000100010",
                            4978 => "100101010",
                            4979 => "110011010",
                            4980 => "011000010",
                            4981 => "101010010",
                            4982 => "011010100",
                            4983 => "100111010",
                            4984 => "100111000",
                            4985 => "111100000",
                            4986 => "000010110",
                            4987 => "001101000",
                            4988 => "001100000",
                            4989 => "100000100",
                            4990 => "010001010",
                            4991 => "100101110",
                            4992 => "010100000",
                            4993 => "000100100",
                            4994 => "110010000",
                            4995 => "111110110",
                            4996 => "001110100",
                            4997 => "111000000",
                            4998 => "001011000",
                            4999 => "001100110",
                            5000 => "100001110",
                            5001 => "101001100",
                            5002 => "110111110",
                            5003 => "001010000",
                            5004 => "100000100",
                            5005 => "011010010",
                            5006 => "110001010",
                            5007 => "000000110",
                            5008 => "111100110",
                            5009 => "111111000",
                            5010 => "000110100",
                            5011 => "001011100",
                            5012 => "010001000",
                            5013 => "011100110",
                            5014 => "100001100",
                            5015 => "110110100",
                            5016 => "111100010",
                            5017 => "100110000",
                            5018 => "111111100",
                            5019 => "010110100",
                            5020 => "000010000",
                            5021 => "011001000",
                            5022 => "010100010",
                            5023 => "111110000",
                            5024 => "011010110",
                            5025 => "100001100",
                            5026 => "111010000",
                            5027 => "000010100",
                            5028 => "100010100",
                            5029 => "000110100",
                            5030 => "101010110",
                            5031 => "001110000",
                            5032 => "110101010",
                            5033 => "100111000",
                            5034 => "011011100",
                            5035 => "001000010",
                            5036 => "001010110",
                            5037 => "001100010",
                            5038 => "010111010",
                            5039 => "101010110",
                            5040 => "101111010",
                            5041 => "000010010",
                            5042 => "100111010",
                            5043 => "111100000",
                            5044 => "010000000",
                            5045 => "010100110",
                            5046 => "111110110",
                            5047 => "111000010",
                            5048 => "110010100",
                            5049 => "001001000",
                            5050 => "000001110",
                            5051 => "101101010",
                            5052 => "010001000",
                            5053 => "011110000",
                            5054 => "011010010",
                            5055 => "111101100",
                            5056 => "101111110",
                            5057 => "110111010",
                            5058 => "110010000",
                            5059 => "000001010",
                            5060 => "111111010",
                            5061 => "101001110",
                            5062 => "001000000",
                            5063 => "111101100",
                            5064 => "111111110",
                            5065 => "011001010",
                            5066 => "000111010",
                            5067 => "100011010",
                            5068 => "011101010",
                            5069 => "111001010",
                            5070 => "011011100",
                            5071 => "101111110",
                            5072 => "101010010",
                            5073 => "101111100",
                            5074 => "110011100",
                            5075 => "010101100",
                            5076 => "011010000",
                            5077 => "111011100",
                            5078 => "101110010",
                            5079 => "000001010",
                            5080 => "010111100",
                            5081 => "111100000",
                            5082 => "111001010",
                            5083 => "100001000",
                            5084 => "101110100",
                            5085 => "000010000",
                            5086 => "001000100",
                            5087 => "111011100",
                            5088 => "101001100",
                            5089 => "010100000",
                            5090 => "101011110",
                            5091 => "000000000",
                            5092 => "111110110",
                            5093 => "100000110",
                            5094 => "101110100",
                            5095 => "011111110",
                            5096 => "110000110",
                            5097 => "001101010",
                            5098 => "011111100",
                            5099 => "100000010",
                            5100 => "011001110",
                            5101 => "100011000",
                            5102 => "000000000",
                            5103 => "011110000",
                            5104 => "001001010",
                            5105 => "111101010",
                            5106 => "101110010",
                            5107 => "011111110",
                            5108 => "101100110",
                            5109 => "000100010",
                            5110 => "000010110",
                            5111 => "111101010",
                            5112 => "101011000",
                            5113 => "011100010",
                            5114 => "000111100",
                            5115 => "001010100",
                            5116 => "011111010",
                            5117 => "111011000",
                            5118 => "010011100",
                            5119 => "000110010",
                            5120 => "110010100",
                            5121 => "100101100",
                            5122 => "110011000",
                            5123 => "111000110",
                            5124 => "000101110",
                            5125 => "011101100",
                            5126 => "101101110",
                            5127 => "111010010",
                            5128 => "010001110",
                            5129 => "001100010",
                            5130 => "110000010",
                            5131 => "011010000",
                            5132 => "110011010",
                            5133 => "010000100",
                            5134 => "001010000",
                            5135 => "101011010",
                            5136 => "010001010",
                            5137 => "100011100",
                            5138 => "011111100",
                            5139 => "000000010",
                            5140 => "000100000",
                            5141 => "010000110",
                            5142 => "101100000",
                            5143 => "110010110",
                            5144 => "001010100",
                            5145 => "000111000",
                            5146 => "111110010",
                            5147 => "000001000",
                            5148 => "011101100",
                            5149 => "100101010",
                            5150 => "111111000",
                            5151 => "000011100",
                            5152 => "100001000",
                            5153 => "110100100",
                            5154 => "000100010",
                            5155 => "011010000",
                            5156 => "101001010",
                            5157 => "010011100",
                            5158 => "011011110",
                            5159 => "000101100",
                            5160 => "000011000",
                            5161 => "011101010",
                            5162 => "011001110",
                            5163 => "111111000",
                            5164 => "110100100",
                            5165 => "001111010",
                            5166 => "000011000",
                            5167 => "010011100",
                            5168 => "001110100",
                            5169 => "011111100",
                            5170 => "010010010",
                            5171 => "100101000",
                            5172 => "110110100",
                            5173 => "010001100",
                            5174 => "000100000",
                            5175 => "000110000",
                            5176 => "110101110",
                            5177 => "110111000",
                            5178 => "010110010",
                            5179 => "101001010",
                            5180 => "100010100",
                            5181 => "001110110",
                            5182 => "000010110",
                            5183 => "101000010",
                            5184 => "110000110",
                            5185 => "011101000",
                            5186 => "111110100",
                            5187 => "011110010",
                            5188 => "111011100",
                            5189 => "111111100",
                            5190 => "001101100",
                            5191 => "010011000",
                            5192 => "111101010",
                            5193 => "101000000",
                            5194 => "110010010",
                            5195 => "011010100",
                            5196 => "010100000",
                            5197 => "010010100",
                            5198 => "100110000",
                            5199 => "011001100",
                            5200 => "000011110",
                            5201 => "110101000",
                            5202 => "011101010",
                            5203 => "111100100",
                            5204 => "101100100",
                            5205 => "111101100",
                            5206 => "011100010",
                            5207 => "000100010",
                            5208 => "001011000",
                            5209 => "101101100",
                            5210 => "100100010",
                            5211 => "011100100",
                            5212 => "100100100",
                            5213 => "111001110",
                            5214 => "010101000",
                            5215 => "000110100",
                            5216 => "011000000",
                            5217 => "111110110",
                            5218 => "101000010",
                            5219 => "000110010",
                            5220 => "110011000",
                            5221 => "110110010",
                            5222 => "001100100",
                            5223 => "111100100",
                            5224 => "100010100",
                            5225 => "111111010",
                            5226 => "101101000",
                            5227 => "101000000",
                            5228 => "100100110",
                            5229 => "110000000",
                            5230 => "111011010",
                            5231 => "010110010",
                            5232 => "001101010",
                            5233 => "111001010",
                            5234 => "011111100",
                            5235 => "001000110",
                            5236 => "101011010",
                            5237 => "110110100",
                            5238 => "101011100",
                            5239 => "110101110",
                            5240 => "111010100",
                            5241 => "000000100",
                            5242 => "110000100",
                            5243 => "110000000",
                            5244 => "010110100",
                            5245 => "111111110",
                            5246 => "100110010",
                            5247 => "111010010",
                            5248 => "001001010",
                            5249 => "110010100",
                            5250 => "000110100",
                            5251 => "101111000",
                            5252 => "000110110",
                            5253 => "111100000",
                            5254 => "001101010",
                            5255 => "101010110",
                            5256 => "100010000",
                            5257 => "001001010",
                            5258 => "100100010",
                            5259 => "001111100",
                            5260 => "111110110",
                            5261 => "110010100",
                            5262 => "000101100",
                            5263 => "111100110",
                            5264 => "111010010",
                            5265 => "110000000",
                            5266 => "100100000",
                            5267 => "110100010",
                            5268 => "010010100",
                            5269 => "000101110",
                            5270 => "001011010",
                            5271 => "000010110",
                            5272 => "000100110",
                            5273 => "011110100",
                            5274 => "111000100",
                            5275 => "000010110",
                            5276 => "010100010",
                            5277 => "100010100",
                            5278 => "000010100",
                            5279 => "100000000",
                            5280 => "111111110",
                            5281 => "011011100",
                            5282 => "101010010",
                            5283 => "000000010",
                            5284 => "010001100",
                            5285 => "100010100",
                            5286 => "110110100",
                            5287 => "110101100",
                            5288 => "111101010",
                            5289 => "110110100",
                            5290 => "100011000",
                            5291 => "000000010",
                            5292 => "101100100",
                            5293 => "110010110",
                            5294 => "010001010",
                            5295 => "100101110",
                            5296 => "000010110",
                            5297 => "010101000",
                            5298 => "111010010",
                            5299 => "010001110",
                            5300 => "110000010",
                            5301 => "100111010",
                            5302 => "011101000",
                            5303 => "111100110",
                            5304 => "100011000",
                            5305 => "110000000",
                            5306 => "001001010",
                            5307 => "101101010",
                            5308 => "011100010",
                            5309 => "011001010",
                            5310 => "101101110",
                            5311 => "110011010",
                            5312 => "110111000",
                            5313 => "100001110",
                            5314 => "010110010",
                            5315 => "011010110",
                            5316 => "000000010",
                            5317 => "101011110",
                            5318 => "100110110",
                            5319 => "111100110",
                            5320 => "011010010",
                            5321 => "010011110",
                            5322 => "011011000",
                            5323 => "111110100",
                            5324 => "001000100",
                            5325 => "010110000",
                            5326 => "010110100",
                            5327 => "110101100",
                            5328 => "011010000",
                            5329 => "000000110",
                            5330 => "001011010",
                            5331 => "100010000",
                            5332 => "100001010",
                            5333 => "010000010",
                            5334 => "000010010",
                            5335 => "111011000",
                            5336 => "111000000",
                            5337 => "001111010",
                            5338 => "111011110",
                            5339 => "100001100",
                            5340 => "110111010",
                            5341 => "111101100",
                            5342 => "011001010",
                            5343 => "000101100",
                            5344 => "101011010",
                            5345 => "110011010",
                            5346 => "001011110",
                            5347 => "000101010",
                            5348 => "100011000",
                            5349 => "111000110",
                            5350 => "100010100",
                            5351 => "110010000",
                            5352 => "000101110",
                            5353 => "000011000",
                            5354 => "101110110",
                            5355 => "110100100",
                            5356 => "000011000",
                            5357 => "100010100",
                            5358 => "111011110",
                            5359 => "110111100",
                            5360 => "100001100",
                            5361 => "110100000",
                            5362 => "011011110",
                            5363 => "010111010",
                            5364 => "011010000",
                            5365 => "101110110",
                            5366 => "000111110",
                            5367 => "101101100",
                            5368 => "110111110",
                            5369 => "110010100",
                            5370 => "011001000",
                            5371 => "000110010",
                            5372 => "100111000",
                            5373 => "001011000",
                            5374 => "011100100",
                            5375 => "101000000",
                            5376 => "110000000",
                            5377 => "011101100",
                            5378 => "001101110",
                            5379 => "000101100",
                            5380 => "100101010",
                            5381 => "001110110",
                            5382 => "110101010",
                            5383 => "011100110",
                            5384 => "010100010",
                            5385 => "111101000",
                            5386 => "001000010",
                            5387 => "110110110",
                            5388 => "000000000",
                            5389 => "000000000",
                            5390 => "000011000",
                            5391 => "100111110",
                            5392 => "111100100",
                            5393 => "010101110",
                            5394 => "100111000",
                            5395 => "101101100",
                            5396 => "110100000",
                            5397 => "000101110",
                            5398 => "010010110",
                            5399 => "000010010",
                            5400 => "000010000",
                            5401 => "000000000",
                            5402 => "010001011",
                            5403 => "000000000",
                            5404 => "000000000",
                            5405 => "001010000",
                            5406 => "011101110",
                            5407 => "111111100",
                            5408 => "010000000",
                            5409 => "000000000",
                            5410 => "100000000",
                            5411 => "000001100",
                            5412 => "101101000",
                            5413 => "010110110",
                            5414 => "000010100",
                            5415 => "110100010",
                            5416 => "111101010",
                            5417 => "011010110",
                            5418 => "010010100",
                            5419 => "011111010",
                            5420 => "100000110",
                            5421 => "101111000",
                            5422 => "111001100",
                            5423 => "101011010",
                            5424 => "000101000",
                            5425 => "011011000",
                            5426 => "110100010",
                            5427 => "010111100",
                            5428 => "111110100",
                            5429 => "010101110",
                            5430 => "011000010",
                            5431 => "010111110",
                            5432 => "011001010",
                            5433 => "100010110",
                            5434 => "010100000",
                            5435 => "000100000",
                            5436 => "000000100",
                            5437 => "000000000",
                            5438 => "010100010",
                            5439 => "101000110",
                            5440 => "000000000",
                            5441 => "000000000",
                            5442 => "100111000",
                            5443 => "101101100",
                            5444 => "110100000",
                            5445 => "000101110",
                            5446 => "010010110",
                            5447 => "000010010",
                            5448 => "000000000",
                            5449 => "001001110",
                            5450 => "100100000",
                            5451 => "111001100",
                            5452 => "001000010",
                            5453 => "010101110",
                            5454 => "000010000",
                            5455 => "000000000",
                            5456 => "010001011",
                            5457 => "000000000",
                            5458 => "000000000",
                            5459 => "011111010",
                            5460 => "110111000",
                            5461 => "010100110",
                            5462 => "010000000",
                            5463 => "000000000",
                            5464 => "001101000",
                            5465 => "000001100",
                            5466 => "001111100",
                            5467 => "011000010",
                            5468 => "101000100",
                            5469 => "100111110",
                            5470 => "100010000",
                            5471 => "111010100",
                            5472 => "000010100",
                            5473 => "110100010",
                            5474 => "111101010",
                            5475 => "011010110",
                            5476 => "000000010",
                            5477 => "101110110",
                            5478 => "111001110",
                            5479 => "000101110",
                            5480 => "000011110",
                            5481 => "001010110",
                            5482 => "100100110",
                            5483 => "101101110",
                            5484 => "011101110",
                            5485 => "001011010",
                            5486 => "101000110",
                            5487 => "110001100",
                            5488 => "010100000",
                            5489 => "000110000",
                            5490 => "000000000",
                            5491 => "010101000",
                            5492 => "111001110",
                            5493 => "011100110",
                            5494 => "000000000",
                            5495 => "000000000",
                            5496 => "000101110",
                            5497 => "000000110",
                            5498 => "000000110",
                            5499 => "000000000",
                            5500 => "010100000",
                            5501 => "001011010",
                            5502 => "101111100",
                            5503 => "111001000",
                            5504 => "110110010",
                            5505 => "000111100",
                            5506 => "111110110",
                            5507 => "101000100",
                            5508 => "111110000",
                            5509 => "010011110",
                            5510 => "100111000",
                            5511 => "011111110",
                            5512 => "100011110",
                            5513 => "101100000",
                            5514 => "011100100",
                            5515 => "001001000",
                            5516 => "111011110",
                            5517 => "000000110",
                            5518 => "110001100",
                            5519 => "000010010",
                            5520 => "010001010",
                            5521 => "101011100",
                            5522 => "111111110",
                            5523 => "011011010",
                            5524 => "001001010",
                            5525 => "100001110",
                            5526 => "100001100",
                            5527 => "000100010",
                            5528 => "000100010",
                            5529 => "100111010",
                            5530 => "100010010",
                            5531 => "111101100",
                            5532 => "110101000",
                            5533 => "010010000",
                            5534 => "101011100",
                            5535 => "101000100",
                            5536 => "110000000",
                            5537 => "011010110",
                            5538 => "111011100",
                            5539 => "111010010",
                            5540 => "101101110",
                            5541 => "011111000",
                            5542 => "011000110",
                            5543 => "110101110",
                            5544 => "101000010",
                            5545 => "011001010",
                            5546 => "100011110",
                            5547 => "101001100",
                            5548 => "110101100",
                            5549 => "101011000",
                            5550 => "011011000",
                            5551 => "110000110",
                            5552 => "100011010",
                            5553 => "110111110",
                            5554 => "011010000",
                            5555 => "001001000",
                            5556 => "100101100",
                            5557 => "110011100",
                            5558 => "111110010",
                            5559 => "101000110",
                            5560 => "101100100",
                            5561 => "101110010",
                            5562 => "101110000",
                            5563 => "000101110",
                            5564 => "100111110",
                            5565 => "110000110",
                            5566 => "111010010",
                            5567 => "101100000",
                            5568 => "000110100",
                            5569 => "000001000",
                            5570 => "010110110",
                            5571 => "111010010",
                            5572 => "110110010",
                            5573 => "110111010",
                            5574 => "100010110",
                            5575 => "010001110",
                            5576 => "111110010",
                            5577 => "000111000",
                            5578 => "111111000",
                            5579 => "011011110",
                            5580 => "000100100",
                            5581 => "000000000",
                            5582 => "000000000",
                            5583 => "000011000",
                            5584 => "100111110",
                            5585 => "111100100",
                            5586 => "010101110",
                            5587 => "100111000",
                            5588 => "101101100",
                            5589 => "110100000",
                            5590 => "000101110",
                            5591 => "010010110",
                            5592 => "000010010",
                            5593 => "000010000",
                            5594 => "000000000",
                            5595 => "010001011",
                            5596 => "000000000",
                            5597 => "000000000",
                            5598 => "001010000",
                            5599 => "100101010",
                            5600 => "001101100",
                            5601 => "010000000",
                            5602 => "000000000",
                            5603 => "100000000",
                            5604 => "000001100",
                            5605 => "001110010",
                            5606 => "110100110",
                            5607 => "000010100",
                            5608 => "110100010",
                            5609 => "111101010",
                            5610 => "011010110",
                            5611 => "101000100",
                            5612 => "100111110",
                            5613 => "100010000",
                            5614 => "111010100",
                            5615 => "111001110",
                            5616 => "000101110",
                            5617 => "000000010",
                            5618 => "101110110",
                            5619 => "011101110",
                            5620 => "001011010",
                            5621 => "101000110",
                            5622 => "110001100",
                            5623 => "000011110",
                            5624 => "001010110",
                            5625 => "100101000",
                            5626 => "000011000",
                            5627 => "010100000",
                            5628 => "000100000",
                            5629 => "000000100",
                            5630 => "000000000",
                            5631 => "110110110",
                            5632 => "000011110",
                            5633 => "000000000",
                            5634 => "000000000",
                            5635 => "000000000",
                            5636 => "000000000",
                            5637 => "000011000",
                            5638 => "100111110",
                            5639 => "111100100",
                            5640 => "010101110",
                            5641 => "100111000",
                            5642 => "101101100",
                            5643 => "110100000",
                            5644 => "000101110",
                            5645 => "010010110",
                            5646 => "000010010",
                            5647 => "000010000",
                            5648 => "000000000",
                            5649 => "010001011",
                            5650 => "100110000",
                            5651 => "000000000",
                            5652 => "010001010",
                            5653 => "111100100",
                            5654 => "011100000",
                            5655 => "010000000",
                            5656 => "000000000",
                            5657 => "100000000",
                            5658 => "000001100",
                            5659 => "101000000",
                            5660 => "010010100",
                            5661 => "000010100",
                            5662 => "110100010",
                            5663 => "111101010",
                            5664 => "011010110",
                            5665 => "000111110",
                            5666 => "000011010",
                            5667 => "010010000",
                            5668 => "000101100",
                            5669 => "111101000",
                            5670 => "000110100",
                            5671 => "000000010",
                            5672 => "101110110",
                            5673 => "111010100",
                            5674 => "000110010",
                            5675 => "110001000",
                            5676 => "101000010",
                            5677 => "111000000",
                            5678 => "111101100",
                            5679 => "000111110",
                            5680 => "010001010",
                            5681 => "010100000",
                            5682 => "000110000",
                            5683 => "000000010",
                            5684 => "111111110",
                            5685 => "101001000",
                            5686 => "000100000",
                            5687 => "000000000",
                            5688 => "000000000",
                            5689 => "000101110",
                            5690 => "000000110",
                            5691 => "000000110",
                            5692 => "000000000",
                            5693 => "000110000",
                            5694 => "000110100",
                            5695 => "011011110",
                            5696 => "010011000",
                            5697 => "111111100",
                            5698 => "111001110",
                            5699 => "100100110",
                            5700 => "101111110",
                            5701 => "010111010",
                            5702 => "001100010",
                            5703 => "100000100",
                            5704 => "011001000",
                            5705 => "110100010",
                            5706 => "000101010",
                            5707 => "111000100",
                            5708 => "001011110",
                            5709 => "110100110",
                            5710 => "111000000",
                            5711 => "101011000",
                            5712 => "100010100",
                            5713 => "000100100",
                            5714 => "011011100",
                            5715 => "000110100",
                            5716 => "101011000",
                            5717 => "100010010",
                            5718 => "000000000",
                            5719 => "000000000",
                            5720 => "000011000",
                            5721 => "100111110",
                            5722 => "111100100",
                            5723 => "010101110",
                            5724 => "100111000",
                            5725 => "101101100",
                            5726 => "110100000",
                            5727 => "000101110",
                            5728 => "010010110",
                            5729 => "000010010",
                            5730 => "000010000",
                            5731 => "000000000",
                            5732 => "010001011",
                            5733 => "100110000",
                            5734 => "000000000",
                            5735 => "010001010",
                            5736 => "111100100",
                            5737 => "011100010",
                            5738 => "010000000",
                            5739 => "000000000",
                            5740 => "100000000",
                            5741 => "000001100",
                            5742 => "101000000",
                            5743 => "010010010",
                            5744 => "000010100",
                            5745 => "110100010",
                            5746 => "111101010",
                            5747 => "011010110",
                            5748 => "000111110",
                            5749 => "000011010",
                            5750 => "010010000",
                            5751 => "000101100",
                            5752 => "111001110",
                            5753 => "000111000",
                            5754 => "000000010",
                            5755 => "101110110",
                            5756 => "101110100",
                            5757 => "101001010",
                            5758 => "100100000",
                            5759 => "110011100",
                            5760 => "010000010",
                            5761 => "110001000",
                            5762 => "010100100",
                            5763 => "000001110",
                            5764 => "010100000",
                            5765 => "000110000",
                            5766 => "000000100",
                            5767 => "000000000",
                            5768 => "110111100",
                            5769 => "110000000",
                            5770 => "000000000",
                            5771 => "000000000",
                            5772 => "000101110",
                            5773 => "000000110",
                            5774 => "000000110",
                            5775 => "000000000",
                            5776 => "000110000",
                            5777 => "100000110",
                            5778 => "001001100",
                            5779 => "101011100",
                            5780 => "000111100",
                            5781 => "010000100",
                            5782 => "011000100",
                            5783 => "101000000",
                            5784 => "110111010",
                            5785 => "100100010",
                            5786 => "000101010",
                            5787 => "000000000",
                            5788 => "001111110",
                            5789 => "010101000",
                            5790 => "011110100",
                            5791 => "101010010",
                            5792 => "000001110",
                            5793 => "010000000",
                            5794 => "010000100",
                            5795 => "010101010",
                            5796 => "011011110",
                            5797 => "011100110",
                            5798 => "001111010",
                            5799 => "110010000",
                            5800 => "001000100",
                            5801 => "100111000",
                            5802 => "101101100",
                            5803 => "110100000",
                            5804 => "000101110",
                            5805 => "010010110",
                            5806 => "000010010",
                            5807 => "000000000",
                            5808 => "001001110",
                            5809 => "100100000",
                            5810 => "111001100",
                            5811 => "001000010",
                            5812 => "010101110",
                            5813 => "000010000",
                            5814 => "000000000",
                            5815 => "010001011",
                            5816 => "000000000",
                            5817 => "000000000",
                            5818 => "001010000",
                            5819 => "110011000",
                            5820 => "011000100",
                            5821 => "010000000",
                            5822 => "000000000",
                            5823 => "010100010",
                            5824 => "000001100",
                            5825 => "111101100",
                            5826 => "000011010",
                            5827 => "000111110",
                            5828 => "000011010",
                            5829 => "010010000",
                            5830 => "000101100",
                            5831 => "000010100",
                            5832 => "110100010",
                            5833 => "111101010",
                            5834 => "011010110",
                            5835 => "000000010",
                            5836 => "101110110",
                            5837 => "111101000",
                            5838 => "000110100",
                            5839 => "111000000",
                            5840 => "111101100",
                            5841 => "000111110",
                            5842 => "010001010",
                            5843 => "111010100",
                            5844 => "000110010",
                            5845 => "110001000",
                            5846 => "101111100",
                            5847 => "010100000",
                            5848 => "000100000",
                            5849 => "000000010",
                            5850 => "001001110",
                            5851 => "101000100",
                            5852 => "011000110",
                            5853 => "000000000",
                            5854 => "000000000",
                            5855 => "100111000",
                            5856 => "101101100",
                            5857 => "110100000",
                            5858 => "000101110",
                            5859 => "010010110",
                            5860 => "000010010",
                            5861 => "000000000",
                            5862 => "001001110",
                            5863 => "100100000",
                            5864 => "111001100",
                            5865 => "001000010",
                            5866 => "010101110",
                            5867 => "000010000",
                            5868 => "000000000",
                            5869 => "010001011",
                            5870 => "000000000",
                            5871 => "000000000",
                            5872 => "001010000",
                            5873 => "100100000",
                            5874 => "011101100",
                            5875 => "010000000",
                            5876 => "000000000",
                            5877 => "010100010",
                            5878 => "000001100",
                            5879 => "001100010",
                            5880 => "111110100",
                            5881 => "000111110",
                            5882 => "000011010",
                            5883 => "010010000",
                            5884 => "000101100",
                            5885 => "000010100",
                            5886 => "110100010",
                            5887 => "111101010",
                            5888 => "011010110",
                            5889 => "000000010",
                            5890 => "101110110",
                            5891 => "111001110",
                            5892 => "000111000",
                            5893 => "010000010",
                            5894 => "110001000",
                            5895 => "010100100",
                            5896 => "000001110",
                            5897 => "101110100",
                            5898 => "101001010",
                            5899 => "100100000",
                            5900 => "111010110",
                            5901 => "010100000",
                            5902 => "000100000",
                            5903 => "000000010",
                            5904 => "001001110",
                            5905 => "011111110",
                            5906 => "000110010",
                            5907 => "000000000",
                            5908 => "000000000",
                            5909 => "100111000",
                            5910 => "101101100",
                            5911 => "110100000",
                            5912 => "000101110",
                            5913 => "010010110",
                            5914 => "000010010",
                            5915 => "000000000",
                            5916 => "001001110",
                            5917 => "100100000",
                            5918 => "111001100",
                            5919 => "001000010",
                            5920 => "010101110",
                            5921 => "000010000",
                            5922 => "000000000",
                            5923 => "010001011",
                            5924 => "000000000",
                            5925 => "000000000",
                            5926 => "010000010",
                            5927 => "110011000",
                            5928 => "011000110",
                            5929 => "010000000",
                            5930 => "000000000",
                            5931 => "010100010",
                            5932 => "000001100",
                            5933 => "111101010",
                            5934 => "111100110",
                            5935 => "000111110",
                            5936 => "000011010",
                            5937 => "010010000",
                            5938 => "000101100",
                            5939 => "000010100",
                            5940 => "110100010",
                            5941 => "111101010",
                            5942 => "011010110",
                            5943 => "000000010",
                            5944 => "101110110",
                            5945 => "111101000",
                            5946 => "000110100",
                            5947 => "111000000",
                            5948 => "111101100",
                            5949 => "000111110",
                            5950 => "010001010",
                            5951 => "111010100",
                            5952 => "000110010",
                            5953 => "110001000",
                            5954 => "101111100",
                            5955 => "010100000",
                            5956 => "000110000",
                            5957 => "000000010",
                            5958 => "001001110",
                            5959 => "001010100",
                            5960 => "001000010",
                            5961 => "000000000",
                            5962 => "000000000",
                            5963 => "000101110",
                            5964 => "000000110",
                            5965 => "000000110",
                            5966 => "000000000",
                            5967 => "000101000",
                            5968 => "011001110",
                            5969 => "011001100",
                            5970 => "111000100",
                            5971 => "000110000",
                            5972 => "011100100",
                            5973 => "010001110",
                            5974 => "100100110",
                            5975 => "101101000",
                            5976 => "110011000",
                            5977 => "100011000",
                            5978 => "111000000",
                            5979 => "001101010",
                            5980 => "001111100",
                            5981 => "110110100",
                            5982 => "100001010",
                            5983 => "011001010",
                            5984 => "001000100",
                            5985 => "000100110",
                            5986 => "001110110",
                            5987 => "100111000",
                            5988 => "101101100",
                            5989 => "110100000",
                            5990 => "000101110",
                            5991 => "010010110",
                            5992 => "000010010",
                            5993 => "000000000",
                            5994 => "001001110",
                            5995 => "100100000",
                            5996 => "111001100",
                            5997 => "001000010",
                            5998 => "010101110",
                            5999 => "000010000",
                            6000 => "000000000",
                            6001 => "010001011",
                            6002 => "000000000",
                            6003 => "000000000",
                            6004 => "010000010",
                            6005 => "100100000",
                            6006 => "011101110",
                            6007 => "010000000",
                            6008 => "000000000",
                            6009 => "010100010",
                            6010 => "000001100",
                            6011 => "001100010",
                            6012 => "111000000",
                            6013 => "000111110",
                            6014 => "000011010",
                            6015 => "010010000",
                            6016 => "000101100",
                            6017 => "000010100",
                            6018 => "110100010",
                            6019 => "111101010",
                            6020 => "011010110",
                            6021 => "000000010",
                            6022 => "101110110",
                            6023 => "111001110",
                            6024 => "000111000",
                            6025 => "010000010",
                            6026 => "110001000",
                            6027 => "010100100",
                            6028 => "000001110",
                            6029 => "101110100",
                            6030 => "101001010",
                            6031 => "100100000",
                            6032 => "111010110",
                            6033 => "010100000",
                            6034 => "000110000",
                            6035 => "000000010",
                            6036 => "001001110",
                            6037 => "101010100",
                            6038 => "001110010",
                            6039 => "000000000",
                            6040 => "000000000",
                            6041 => "000101110",
                            6042 => "000000110",
                            6043 => "000000110",
                            6044 => "000000000",
                            6045 => "000101000",
                            6046 => "111111100",
                            6047 => "010010100",
                            6048 => "111011000",
                            6049 => "011101110",
                            6050 => "011000110",
                            6051 => "111100110",
                            6052 => "011110110",
                            6053 => "110011100",
                            6054 => "101010010",
                            6055 => "000000100",
                            6056 => "110110010",
                            6057 => "101111010",
                            6058 => "011001100",
                            6059 => "001101010",
                            6060 => "101011110",
                            6061 => "000000110",
                            6062 => "011100000",
                            6063 => "100101100",
                            6064 => "111010000",
                            6065 => "000000000",
                            6066 => "000000000",
                            6067 => "000011000",
                            6068 => "100111110",
                            6069 => "111100100",
                            6070 => "010101110",
                            6071 => "100111000",
                            6072 => "101101100",
                            6073 => "110100000",
                            6074 => "000101110",
                            6075 => "010010110",
                            6076 => "000010010",
                            6077 => "000010000",
                            6078 => "000000000",
                            6079 => "010001011",
                            6080 => "000000000",
                            6081 => "000000000",
                            6082 => "001010000",
                            6083 => "111100100",
                            6084 => "011100100",
                            6085 => "010000000",
                            6086 => "000000000",
                            6087 => "100000000",
                            6088 => "000001100",
                            6089 => "101000000",
                            6090 => "111111010",
                            6091 => "000010100",
                            6092 => "110100010",
                            6093 => "111101010",
                            6094 => "011010110",
                            6095 => "000111110",
                            6096 => "000011010",
                            6097 => "010010000",
                            6098 => "000101100",
                            6099 => "111101000",
                            6100 => "000110100",
                            6101 => "000000010",
                            6102 => "101110110",
                            6103 => "111010100",
                            6104 => "000110010",
                            6105 => "110001000",
                            6106 => "101111100",
                            6107 => "111000000",
                            6108 => "111101100",
                            6109 => "000111110",
                            6110 => "010111100",
                            6111 => "010100000",
                            6112 => "000100000",
                            6113 => "000000010",
                            6114 => "111111110",
                            6115 => "101000010",
                            6116 => "011100100",
                            6117 => "000000000",
                            6118 => "000000000",
                            6119 => "000000000",
                            6120 => "000000000",
                            6121 => "000011000",
                            6122 => "100111110",
                            6123 => "111100100",
                            6124 => "010101110",
                            6125 => "100111000",
                            6126 => "101101100",
                            6127 => "110100000",
                            6128 => "000101110",
                            6129 => "010010110",
                            6130 => "000010010",
                            6131 => "000010000",
                            6132 => "000000000",
                            6133 => "010001011",
                            6134 => "000000000",
                            6135 => "000000000",
                            6136 => "001010000",
                            6137 => "111100100",
                            6138 => "011100110",
                            6139 => "010000000",
                            6140 => "000000000",
                            6141 => "100000000",
                            6142 => "000001100",
                            6143 => "101000000",
                            6144 => "111111000",
                            6145 => "000010100",
                            6146 => "110100010",
                            6147 => "111101010",
                            6148 => "011010110",
                            6149 => "000111110",
                            6150 => "000011010",
                            6151 => "010010000",
                            6152 => "000101100",
                            6153 => "111001110",
                            6154 => "000111000",
                            6155 => "000000010",
                            6156 => "101110110",
                            6157 => "101110100",
                            6158 => "101001010",
                            6159 => "100100000",
                            6160 => "111010110",
                            6161 => "010000010",
                            6162 => "110001000",
                            6163 => "010100100",
                            6164 => "001000000",
                            6165 => "010100000",
                            6166 => "000100000",
                            6167 => "000000100",
                            6168 => "000000000",
                            6169 => "011111100",
                            6170 => "001001110",
                            6171 => "000000000",
                            6172 => "000000000",
                            6173 => "100111000",
                            6174 => "101101100",
                            6175 => "110100000",
                            6176 => "000101110",
                            6177 => "010010110",
                            6178 => "000010010",
                            6179 => "000000000",
                            6180 => "001001110",
                            6181 => "100100000",
                            6182 => "111001100",
                            6183 => "001000010",
                            6184 => "010101110",
                            6185 => "000010000",
                            6186 => "000000000",
                            6187 => "010001011",
                            6188 => "000000000",
                            6189 => "000000000",
                            6190 => "011110000",
                            6191 => "110111000",
                            6192 => "010101000",
                            6193 => "010000000",
                            6194 => "000000000",
                            6195 => "001101000",
                            6196 => "000001100",
                            6197 => "001111100",
                            6198 => "011001010",
                            6199 => "101000100",
                            6200 => "100111110",
                            6201 => "100010000",
                            6202 => "111010100",
                            6203 => "000010100",
                            6204 => "110100010",
                            6205 => "111101010",
                            6206 => "011010110",
                            6207 => "000000010",
                            6208 => "101110110",
                            6209 => "111001110",
                            6210 => "000101110",
                            6211 => "000011110",
                            6212 => "001010110",
                            6213 => "100101000",
                            6214 => "000011000",
                            6215 => "011101110",
                            6216 => "001011010",
                            6217 => "101000110",
                            6218 => "110001100",
                            6219 => "010100000",
                            6220 => "000110000",
                            6221 => "000000000",
                            6222 => "010101000",
                            6223 => "101101110",
                            6224 => "000000000",
                            6225 => "000000000",
                            6226 => "000000000",
                            6227 => "000101110",
                            6228 => "000000110",
                            6229 => "000000110",
                            6230 => "000000000",
                            6231 => "010010110",
                            6232 => "001110100",
                            6233 => "111111010",
                            6234 => "010001100",
                            6235 => "111000100",
                            6236 => "001110110",
                            6237 => "011011100",
                            6238 => "001001100",
                            6239 => "111001100",
                            6240 => "110010100",
                            6241 => "100101010",
                            6242 => "010010000",
                            6243 => "110000100",
                            6244 => "011111010",
                            6245 => "011111110",
                            6246 => "100101100",
                            6247 => "010000000",
                            6248 => "011111000",
                            6249 => "000000100",
                            6250 => "111101000",
                            6251 => "001000100",
                            6252 => "001011110",
                            6253 => "110010110",
                            6254 => "110110110",
                            6255 => "011011000",
                            6256 => "101101100",
                            6257 => "001111100",
                            6258 => "101011100",
                            6259 => "001011000",
                            6260 => "000100110",
                            6261 => "010111110",
                            6262 => "111011110",
                            6263 => "111011100",
                            6264 => "001001010",
                            6265 => "110110000",
                            6266 => "010111000",
                            6267 => "001101000",
                            6268 => "101010100",
                            6269 => "000111100",
                            6270 => "011011000",
                            6271 => "001011110",
                            6272 => "001101110",
                            6273 => "100011110",
                            6274 => "010011100",
                            6275 => "101110010",
                            6276 => "111010010",
                            6277 => "100100110",
                            6278 => "001111100",
                            6279 => "100110000",
                            6280 => "101110010",
                            6281 => "100101110",
                            6282 => "010000110",
                            6283 => "001010100",
                            6284 => "011010010",
                            6285 => "000110110",
                            6286 => "001001010",
                            6287 => "101110110",
                            6288 => "100000010",
                            6289 => "011001100",
                            6290 => "000101110",
                            6291 => "101111010",
                            6292 => "100011010",
                            6293 => "011111110",
                            6294 => "100110100",
                            6295 => "111001100",
                            6296 => "011000100",
                            6297 => "101110100",
                            6298 => "100110100",
                            6299 => "001101000",
                            6300 => "101101100",
                            6301 => "011001000",
                            6302 => "001101100",
                            6303 => "010100000",
                            6304 => "111111010",
                            6305 => "110001100",
                            6306 => "111101100",
                            6307 => "000000000",
                            6308 => "000000000",
                            6309 => "000011000",
                            6310 => "100111110",
                            6311 => "111100100",
                            6312 => "010101110",
                            6313 => "100111000",
                            6314 => "101101100",
                            6315 => "110100000",
                            6316 => "000101110",
                            6317 => "010010110",
                            6318 => "000010010",
                            6319 => "000010000",
                            6320 => "000000000",
                            6321 => "010001011",
                            6322 => "000000000",
                            6323 => "000000000",
                            6324 => "001010000",
                            6325 => "100101010",
                            6326 => "001101110",
                            6327 => "010000000",
                            6328 => "000000000",
                            6329 => "100000000",
                            6330 => "000001100",
                            6331 => "001110010",
                            6332 => "110100100",
                            6333 => "000010100",
                            6334 => "110100010",
                            6335 => "111101010",
                            6336 => "011010110",
                            6337 => "101000100",
                            6338 => "100111110",
                            6339 => "100010000",
                            6340 => "111010100",
                            6341 => "111001110",
                            6342 => "000101110",
                            6343 => "000000010",
                            6344 => "101110110",
                            6345 => "011101110",
                            6346 => "001011010",
                            6347 => "101000110",
                            6348 => "110001100",
                            6349 => "000011110",
                            6350 => "001010110",
                            6351 => "100101000",
                            6352 => "010111000",
                            6353 => "010100000",
                            6354 => "000100000",
                            6355 => "000000010",
                            6356 => "111111110",
                            6357 => "110110100",
                            6358 => "110000000",
                            6359 => "000000000",
                            6360 => "000000000",
                            6361 => "100111000",
                            6362 => "101101100",
                            6363 => "110100000",
                            6364 => "000101110",
                            6365 => "010010110",
                            6366 => "000010010",
                            6367 => "000000000",
                            6368 => "001001110",
                            6369 => "100100000",
                            6370 => "111001100",
                            6371 => "001000010",
                            6372 => "010101110",
                            6373 => "000010000",
                            6374 => "000000000",
                            6375 => "010001011",
                            6376 => "000000000",
                            6377 => "000000000",
                            6378 => "101010000",
                            6379 => "110111000",
                            6380 => "010101010",
                            6381 => "010000000",
                            6382 => "000000000",
                            6383 => "001101000",
                            6384 => "000001100",
                            6385 => "001111100",
                            6386 => "001101000",
                            6387 => "101000100",
                            6388 => "100111110",
                            6389 => "100010000",
                            6390 => "111010100",
                            6391 => "000010100",
                            6392 => "110100010",
                            6393 => "111101010",
                            6394 => "011010110",
                            6395 => "000000010",
                            6396 => "101110110",
                            6397 => "111001110",
                            6398 => "000101110",
                            6399 => "000011110",
                            6400 => "001010110",
                            6401 => "100101000",
                            6402 => "010111000",
                            6403 => "011101110",
                            6404 => "001011010",
                            6405 => "101000110",
                            6406 => "110001100",
                            6407 => "010100000",
                            6408 => "000110000",
                            6409 => "000000000",
                            6410 => "010101000",
                            6411 => "111001100",
                            6412 => "001000100",
                            6413 => "000000000",
                            6414 => "000000000",
                            6415 => "000101110",
                            6416 => "000000110",
                            6417 => "000000110",
                            6418 => "000000000",
                            6419 => "011110110",
                            6420 => "101101010",
                            6421 => "001111000",
                            6422 => "100110010",
                            6423 => "110000000",
                            6424 => "100001110",
                            6425 => "101000110",
                            6426 => "110011110",
                            6427 => "011100010",
                            6428 => "010000100",
                            6429 => "010001100",
                            6430 => "100000010",
                            6431 => "100010110",
                            6432 => "101101010",
                            6433 => "111110000",
                            6434 => "101101100",
                            6435 => "000011110",
                            6436 => "010100000",
                            6437 => "110111100",
                            6438 => "011011100",
                            6439 => "110011100",
                            6440 => "101110110",
                            6441 => "101011110",
                            6442 => "111000110",
                            6443 => "110000110",
                            6444 => "011011100",
                            6445 => "010010010",
                            6446 => "111101000",
                            6447 => "110111000",
                            6448 => "101000110",
                            6449 => "101101000",
                            6450 => "000000010",
                            6451 => "111010100",
                            6452 => "101000010",
                            6453 => "101110110",
                            6454 => "011010010",
                            6455 => "011101110",
                            6456 => "110001000",
                            6457 => "100010010",
                            6458 => "001011110",
                            6459 => "101000110",
                            6460 => "111111110",
                            6461 => "001100010",
                            6462 => "101100100",
                            6463 => "000010010",
                            6464 => "100000110",
                            6465 => "101100000",
                            6466 => "100110100",
                            6467 => "000001100",
                            6468 => "101011110",
                            6469 => "101111000",
                            6470 => "101111010",
                            6471 => "100110000",
                            6472 => "101111000",
                            6473 => "000111000",
                            6474 => "001100110",
                            6475 => "010000100",
                            6476 => "001011100",
                            6477 => "001011010",
                            6478 => "111000000",
                            6479 => "011010100",
                            6480 => "110110000",
                            6481 => "100000110",
                            6482 => "111000100",
                            6483 => "100101010",
                            6484 => "010001110",
                            6485 => "011010010",
                            6486 => "000111110",
                            6487 => "110110100",
                            6488 => "101110000",
                            6489 => "000001000",
                            6490 => "110101100",
                            6491 => "110001110",
                            6492 => "101110000",
                            6493 => "100011100",
                            6494 => "110100010",
                            6495 => "101111100",
                            6496 => "011110100",
                            6497 => "011110100",
                            6498 => "110000100",
                            6499 => "110010110",
                            6500 => "101010000",
                            6501 => "001110100",
                            6502 => "000000110",
                            6503 => "111111110",
                            6504 => "011100100",
                            6505 => "000010100",
                            6506 => "111111010",
                            6507 => "110110100",
                            6508 => "100110110",
                            6509 => "010011110",
                            6510 => "101001100",
                            6511 => "011100000",
                            6512 => "101110000",
                            6513 => "000111010",
                            6514 => "101110010",
                            6515 => "101001100",
                            6516 => "001000010",
                            6517 => "010000000",
                            6518 => "111000100",
                            6519 => "011000000",
                            6520 => "011111100",
                            6521 => "011011110",
                            6522 => "000011010",
                            6523 => "110100110",
                            6524 => "101000100",
                            6525 => "010000110",
                            6526 => "100010100",
                            6527 => "011010110",
                            6528 => "010011010",
                            6529 => "011110000",
                            6530 => "001000110",
                            6531 => "010101110",
                            6532 => "000000000",
                            6533 => "100111100",
                            6534 => "000111000",
                            6535 => "110110010",
                            6536 => "101100100",
                            6537 => "101101100",
                            6538 => "011100000",
                            6539 => "110101010",
                            6540 => "101100000",
                            6541 => "001001110",
                            6542 => "110111110",
                            6543 => "000000000",
                            6544 => "000000000",
                            6545 => "000011000",
                            6546 => "100111110",
                            6547 => "111100100",
                            6548 => "010101110",
                            6549 => "100111000",
                            6550 => "101101100",
                            6551 => "110100000",
                            6552 => "000101110",
                            6553 => "010010110",
                            6554 => "000010010",
                            6555 => "000010000",
                            6556 => "000000000",
                            6557 => "010001011",
                            6558 => "000000000",
                            6559 => "000000000",
                            6560 => "001010000",
                            6561 => "100101010",
                            6562 => "001110000",
                            6563 => "010000000",
                            6564 => "000000000",
                            6565 => "100000000",
                            6566 => "000001100",
                            6567 => "001110010",
                            6568 => "110100010",
                            6569 => "000010100",
                            6570 => "110100010",
                            6571 => "111101010",
                            6572 => "011010110",
                            6573 => "101000100",
                            6574 => "100111110",
                            6575 => "100010000",
                            6576 => "111010100",
                            6577 => "111001110",
                            6578 => "000101110",
                            6579 => "000000010",
                            6580 => "101110110",
                            6581 => "011101110",
                            6582 => "001011010",
                            6583 => "101000110",
                            6584 => "110001100",
                            6585 => "000011110",
                            6586 => "001010110",
                            6587 => "100101000",
                            6588 => "110111000",
                            6589 => "010100000",
                            6590 => "000100000",
                            6591 => "000000010",
                            6592 => "111111110",
                            6593 => "110110100",
                            6594 => "010000000",
                            6595 => "000000000",
                            6596 => "000000000",
                            6597 => "100111000",
                            6598 => "101101100",
                            6599 => "110100000",
                            6600 => "000101110",
                            6601 => "010010110",
                            6602 => "000010010",
                            6603 => "000000000",
                            6604 => "001001110",
                            6605 => "100100000",
                            6606 => "111001100",
                            6607 => "001000010",
                            6608 => "010101110",
                            6609 => "000010000",
                            6610 => "000000000",
                            6611 => "010001011",
                            6612 => "000000000",
                            6613 => "000000000",
                            6614 => "100101110",
                            6615 => "110111000",
                            6616 => "010101100",
                            6617 => "010000000",
                            6618 => "000000000",
                            6619 => "001101000",
                            6620 => "000001100",
                            6621 => "001111100",
                            6622 => "010001000",
                            6623 => "101000100",
                            6624 => "100111110",
                            6625 => "100010000",
                            6626 => "111010100",
                            6627 => "000010100",
                            6628 => "110100010",
                            6629 => "111101010",
                            6630 => "011010110",
                            6631 => "000000010",
                            6632 => "101110110",
                            6633 => "111001110",
                            6634 => "000101110",
                            6635 => "000011110",
                            6636 => "001010110",
                            6637 => "100101000",
                            6638 => "110111000",
                            6639 => "011101110",
                            6640 => "001011010",
                            6641 => "101000110",
                            6642 => "110001100",
                            6643 => "010100000",
                            6644 => "000110000",
                            6645 => "000000000",
                            6646 => "010101000",
                            6647 => "101111110",
                            6648 => "010111110",
                            6649 => "000000000",
                            6650 => "000000000",
                            6651 => "000101110",
                            6652 => "000000110",
                            6653 => "000000110",
                            6654 => "000000000",
                            6655 => "011010100",
                            6656 => "001010010",
                            6657 => "110000010",
                            6658 => "000011010",
                            6659 => "011100000",
                            6660 => "100010100",
                            6661 => "010110010",
                            6662 => "011001000",
                            6663 => "110110010",
                            6664 => "110010000",
                            6665 => "101010100",
                            6666 => "100100100",
                            6667 => "000011010",
                            6668 => "001101110",
                            6669 => "010100100",
                            6670 => "100100010",
                            6671 => "110010010",
                            6672 => "011110110",
                            6673 => "101110000",
                            6674 => "000011000",
                            6675 => "101111100",
                            6676 => "011010100",
                            6677 => "001100100",
                            6678 => "110101110",
                            6679 => "001100010",
                            6680 => "011101000",
                            6681 => "110111010",
                            6682 => "000011000",
                            6683 => "010000100",
                            6684 => "000011000",
                            6685 => "101000010",
                            6686 => "101011010",
                            6687 => "000110110",
                            6688 => "101110010",
                            6689 => "000101110",
                            6690 => "011110010",
                            6691 => "001110010",
                            6692 => "000101110",
                            6693 => "010001110",
                            6694 => "100110100",
                            6695 => "101001110",
                            6696 => "001011100",
                            6697 => "110010010",
                            6698 => "010110100",
                            6699 => "000010000",
                            6700 => "111011010",
                            6701 => "000111010",
                            6702 => "000110100",
                            6703 => "100010010",
                            6704 => "010111010",
                            6705 => "111000010",
                            6706 => "000101010",
                            6707 => "000111010",
                            6708 => "000000100",
                            6709 => "000110000",
                            6710 => "111111100",
                            6711 => "001011010",
                            6712 => "100001000",
                            6713 => "101011010",
                            6714 => "011100000",
                            6715 => "011011110",
                            6716 => "010100000",
                            6717 => "101100000",
                            6718 => "100001100",
                            6719 => "001011100",
                            6720 => "000001010",
                            6721 => "101101100",
                            6722 => "000101100",
                            6723 => "010111100",
                            6724 => "001000100",
                            6725 => "100101010",
                            6726 => "001110000",
                            6727 => "101000100",
                            6728 => "011010110",
                            6729 => "111000110",
                            6730 => "011101100",
                            6731 => "111000010",
                            6732 => "100001000",
                            6733 => "100000110",
                            6734 => "001010100",
                            6735 => "100001010",
                            6736 => "110111000",
                            6737 => "100011010",
                            6738 => "010001010",
                            6739 => "101110100",
                            6740 => "010101100",
                            6741 => "000100010",
                            6742 => "001001110",
                            6743 => "000100100",
                            6744 => "010101100",
                            6745 => "111000110",
                            6746 => "101111010",
                            6747 => "111001010",
                            6748 => "000000010",
                            6749 => "110011000",
                            6750 => "100101110",
                            6751 => "010000100",
                            6752 => "110010010",
                            6753 => "000111100",
                            6754 => "101000010",
                            6755 => "111001110",
                            6756 => "000000010",
                            6757 => "011001100",
                            6758 => "010001000",
                            6759 => "101000110",
                            6760 => "000001110",
                            6761 => "010001000",
                            6762 => "000000000",
                            6763 => "000000000",
                            6764 => "000011000",
                            6765 => "100111110",
                            6766 => "111100100",
                            6767 => "010101110",
                            6768 => "100111000",
                            6769 => "101101100",
                            6770 => "110100000",
                            6771 => "000101110",
                            6772 => "010010110",
                            6773 => "000010010",
                            6774 => "000010000",
                            6775 => "000000000",
                            6776 => "010001011",
                            6777 => "000000000",
                            6778 => "000000000",
                            6779 => "001010000",
                            6780 => "100101010",
                            6781 => "001110010",
                            6782 => "010000000",
                            6783 => "000000000",
                            6784 => "100000000",
                            6785 => "000001100",
                            6786 => "001110010",
                            6787 => "110100000",
                            6788 => "000010100",
                            6789 => "110100010",
                            6790 => "111101010",
                            6791 => "011010110",
                            6792 => "101000100",
                            6793 => "100111110",
                            6794 => "100010000",
                            6795 => "111010100",
                            6796 => "111001110",
                            6797 => "000101110",
                            6798 => "000000010",
                            6799 => "101110110",
                            6800 => "011101110",
                            6801 => "001011010",
                            6802 => "101000110",
                            6803 => "110001100",
                            6804 => "000011110",
                            6805 => "001010110",
                            6806 => "100101010",
                            6807 => "010010110",
                            6808 => "010100000",
                            6809 => "000100000",
                            6810 => "000000010",
                            6811 => "111111100",
                            6812 => "110110010",
                            6813 => "110100100",
                            6814 => "000000000",
                            6815 => "000000000",
                            6816 => "000000000",
                            6817 => "000000000",
                            6818 => "000011000",
                            6819 => "100111110",
                            6820 => "111100100",
                            6821 => "010101110",
                            6822 => "100111000",
                            6823 => "101101100",
                            6824 => "110100000",
                            6825 => "000101110",
                            6826 => "010010110",
                            6827 => "000010010",
                            6828 => "000010000",
                            6829 => "000000000",
                            6830 => "010001011",
                            6831 => "100110000",
                            6832 => "000000000",
                            6833 => "010010000",
                            6834 => "111010000",
                            6835 => "001000100",
                            6836 => "010000000",
                            6837 => "000000000",
                            6838 => "100000000",
                            6839 => "000001100",
                            6840 => "101010100",
                            6841 => "101000110",
                            6842 => "000010100",
                            6843 => "110100010",
                            6844 => "111101010",
                            6845 => "011010110",
                            6846 => "000111110",
                            6847 => "000011010",
                            6848 => "010010000",
                            6849 => "000010000",
                            6850 => "111101000",
                            6851 => "000110110",
                            6852 => "000000010",
                            6853 => "101110110",
                            6854 => "011000010",
                            6855 => "011110100",
                            6856 => "100000010",
                            6857 => "001110110",
                            6858 => "001000010",
                            6859 => "011111010",
                            6860 => "011011100",
                            6861 => "000100100",
                            6862 => "010100000",
                            6863 => "000110000",
                            6864 => "000000010",
                            6865 => "111111000",
                            6866 => "110111110",
                            6867 => "101001100",
                            6868 => "000000000",
                            6869 => "000000000",
                            6870 => "000101110",
                            6871 => "000000110",
                            6872 => "000000110",
                            6873 => "000000000",
                            6874 => "000110110",
                            6875 => "000110010",
                            6876 => "011000100",
                            6877 => "110011110",
                            6878 => "110111100",
                            6879 => "010011100",
                            6880 => "001001000",
                            6881 => "101010000",
                            6882 => "100111000",
                            6883 => "010101000",
                            6884 => "111000010",
                            6885 => "111001010",
                            6886 => "110101000",
                            6887 => "101111100",
                            6888 => "111000000",
                            6889 => "111111100",
                            6890 => "011011000",
                            6891 => "000110100",
                            6892 => "011111110",
                            6893 => "100101100",
                            6894 => "011110100",
                            6895 => "111000100",
                            6896 => "111001000",
                            6897 => "100101010",
                            6898 => "110101110",
                            6899 => "101010010",
                            6900 => "000011000",
                            6901 => "111011100",
                            6902 => "100111000",
                            6903 => "101101100",
                            6904 => "110100000",
                            6905 => "000101110",
                            6906 => "010010110",
                            6907 => "000010010",
                            6908 => "000000000",
                            6909 => "001001110",
                            6910 => "100100000",
                            6911 => "111001100",
                            6912 => "001000010",
                            6913 => "010101110",
                            6914 => "000010000",
                            6915 => "000000000",
                            6916 => "010001011",
                            6917 => "000000000",
                            6918 => "000000010",
                            6919 => "010011000",
                            6920 => "110111000",
                            6921 => "010101110",
                            6922 => "010000000",
                            6923 => "000000000",
                            6924 => "001101000",
                            6925 => "000001100",
                            6926 => "001111010",
                            6927 => "100011100",
                            6928 => "101000100",
                            6929 => "100111110",
                            6930 => "100010000",
                            6931 => "111010100",
                            6932 => "000010100",
                            6933 => "110100010",
                            6934 => "111101010",
                            6935 => "011010110",
                            6936 => "000000010",
                            6937 => "101110110",
                            6938 => "111001110",
                            6939 => "000101110",
                            6940 => "000011110",
                            6941 => "001010110",
                            6942 => "100101010",
                            6943 => "010010110",
                            6944 => "011101110",
                            6945 => "001011010",
                            6946 => "101000110",
                            6947 => "110001100",
                            6948 => "010100000",
                            6949 => "000110000",
                            6950 => "000000000",
                            6951 => "010101000",
                            6952 => "100100100",
                            6953 => "011010100",
                            6954 => "000000000",
                            6955 => "000000000",
                            6956 => "000101110",
                            6957 => "000000110",
                            6958 => "000000110",
                            6959 => "000000010",
                            6960 => "000111110",
                            6961 => "011100010",
                            6962 => "110110000",
                            6963 => "001111100",
                            6964 => "011111100",
                            6965 => "001100000",
                            6966 => "000000100",
                            6967 => "111110110",
                            6968 => "111100100",
                            6969 => "010101100",
                            6970 => "001000010",
                            6971 => "110000100",
                            6972 => "000001110",
                            6973 => "111011110",
                            6974 => "010011100",
                            6975 => "000000100",
                            6976 => "001000010",
                            6977 => "010111110",
                            6978 => "001001110",
                            6979 => "110110100",
                            6980 => "110001110",
                            6981 => "101000010",
                            6982 => "100111100",
                            6983 => "000011100",
                            6984 => "100101010",
                            6985 => "011110000",
                            6986 => "110111100",
                            6987 => "100000110",
                            6988 => "101101000",
                            6989 => "000101110",
                            6990 => "100111000",
                            6991 => "000111000",
                            6992 => "000100010",
                            6993 => "101110110",
                            6994 => "001011010",
                            6995 => "001100000",
                            6996 => "011101100",
                            6997 => "001110110",
                            6998 => "000101000",
                            6999 => "111101110",
                            7000 => "101011000",
                            7001 => "011101110",
                            7002 => "111100000",
                            7003 => "110001110",
                            7004 => "110001100",
                            7005 => "110000010",
                            7006 => "011100010",
                            7007 => "101101000",
                            7008 => "111100110",
                            7009 => "010100000",
                            7010 => "000001100",
                            7011 => "011000100",
                            7012 => "010001000",
                            7013 => "101111010",
                            7014 => "011000010",
                            7015 => "111111100",
                            7016 => "010111100",
                            7017 => "011111110",
                            7018 => "011001000",
                            7019 => "001101110",
                            7020 => "001000010",
                            7021 => "000001010",
                            7022 => "100100010",
                            7023 => "011000100",
                            7024 => "110010000",
                            7025 => "111010100",
                            7026 => "110110000",
                            7027 => "001110010",
                            7028 => "000000100",
                            7029 => "111011000",
                            7030 => "110010000",
                            7031 => "110101100",
                            7032 => "111111010",
                            7033 => "010011110",
                            7034 => "100001110",
                            7035 => "000011110",
                            7036 => "111001010",
                            7037 => "101010100",
                            7038 => "110000000",
                            7039 => "110000000",
                            7040 => "111000000",
                            7041 => "000101110",
                            7042 => "100000100",
                            7043 => "000110010",
                            7044 => "111101100",
                            7045 => "001001100",
                            7046 => "111001110",
                            7047 => "010101110",
                            7048 => "011110110",
                            7049 => "010101010",
                            7050 => "001100000",
                            7051 => "111010110",
                            7052 => "001110100",
                            7053 => "100110000",
                            7054 => "101101010",
                            7055 => "101000110",
                            7056 => "100010110",
                            7057 => "101010110",
                            7058 => "100110110",
                            7059 => "010101000",
                            7060 => "101110010",
                            7061 => "000110000",
                            7062 => "111110110",
                            7063 => "010000010",
                            7064 => "000000110",
                            7065 => "111110010",
                            7066 => "011111000",
                            7067 => "100101000",
                            7068 => "101101100",
                            7069 => "100000100",
                            7070 => "001101000",
                            7071 => "111110000",
                            7072 => "001101010",
                            7073 => "010000010",
                            7074 => "011010100",
                            7075 => "100111110",
                            7076 => "000110000",
                            7077 => "101011010",
                            7078 => "101000100",
                            7079 => "100000110",
                            7080 => "101111100",
                            7081 => "011100000",
                            7082 => "010100100",
                            7083 => "010000100",
                            7084 => "001010110",
                            7085 => "111011110",
                            7086 => "111111110",
                            7087 => "001000110",
                            7088 => "000011100",
                            7089 => "010100010",
                            7090 => "011100000",
                            7091 => "001011100",
                            7092 => "010011010",
                            7093 => "111000010",
                            7094 => "000110010",
                            7095 => "110101000",
                            7096 => "100010000",
                            7097 => "010101010",
                            7098 => "100110010",
                            7099 => "001100100",
                            7100 => "111110000",
                            7101 => "100010000",
                            7102 => "111010000",
                            7103 => "100001100",
                            7104 => "110111010",
                            7105 => "100110100",
                            7106 => "011011000",
                            7107 => "001111010",
                            7108 => "010101000",
                            7109 => "011000000",
                            7110 => "110101000",
                            7111 => "111011000",
                            7112 => "111011100",
                            7113 => "111101010",
                            7114 => "110001110",
                            7115 => "000011010",
                            7116 => "111011100",
                            7117 => "100011110",
                            7118 => "111100000",
                            7119 => "111100010",
                            7120 => "100001110",
                            7121 => "111110000",
                            7122 => "110111000",
                            7123 => "001010110",
                            7124 => "000010000",
                            7125 => "010001100",
                            7126 => "010111010",
                            7127 => "101101110",
                            7128 => "001101000",
                            7129 => "101000110",
                            7130 => "011101100",
                            7131 => "101110100",
                            7132 => "111010000",
                            7133 => "101011100",
                            7134 => "001000000",
                            7135 => "010110000",
                            7136 => "101100000",
                            7137 => "011110000",
                            7138 => "100001000",
                            7139 => "011111110",
                            7140 => "000010100",
                            7141 => "010100100",
                            7142 => "010011110",
                            7143 => "100100110",
                            7144 => "000111100",
                            7145 => "101000000",
                            7146 => "110111110",
                            7147 => "001110000",
                            7148 => "100011000",
                            7149 => "101011110",
                            7150 => "100111110",
                            7151 => "111100110",
                            7152 => "101100110",
                            7153 => "101001000",
                            7154 => "011111000",
                            7155 => "011101010",
                            7156 => "001110000",
                            7157 => "100011000",
                            7158 => "100101000",
                            7159 => "111010000",
                            7160 => "110111010",
                            7161 => "011001000",
                            7162 => "100001110",
                            7163 => "001011100",
                            7164 => "110101100",
                            7165 => "011100110",
                            7166 => "011111010",
                            7167 => "111100000",
                            7168 => "110001010",
                            7169 => "110110000",
                            7170 => "101110010",
                            7171 => "110011000",
                            7172 => "000110000",
                            7173 => "110001010",
                            7174 => "000110010",
                            7175 => "111111110",
                            7176 => "001011000",
                            7177 => "011110100",
                            7178 => "111010110",
                            7179 => "010001000",
                            7180 => "100001000",
                            7181 => "001011100",
                            7182 => "101110100",
                            7183 => "101010100",
                            7184 => "001000000",
                            7185 => "001000100",
                            7186 => "100011000",
                            7187 => "100100000",
                            7188 => "100111110",
                            7189 => "010001010",
                            7190 => "001011110",
                            7191 => "111001100",
                            7192 => "011010100",
                            7193 => "000100110",
                            7194 => "110011000",
                            7195 => "111110100",
                            7196 => "000101010",
                            7197 => "110111110",
                            7198 => "011111000",
                            7199 => "101110100",
                            7200 => "101000010",
                            7201 => "011101110",
                            7202 => "000011110",
                            7203 => "000010010",
                            7204 => "111000000",
                            7205 => "010000000",
                            7206 => "001111110",
                            7207 => "011010100",
                            7208 => "100110000",
                            7209 => "000100010",
                            7210 => "110010000",
                            7211 => "011110110",
                            7212 => "010100000",
                            7213 => "000111110",
                            7214 => "100011110",
                            7215 => "001001110",
                            7216 => "110011100",
                            7217 => "000011100",
                            7218 => "000001100",
                            7219 => "000010100",
                            7220 => "101010110",
                            7221 => "011110010",
                            7222 => "101101100",
                            7223 => "101101110",
                            7224 => "010101100",
                            7225 => "111011110",
                            7226 => "101010110",
                            7227 => "110010100",
                            7228 => "001011110",
                            7229 => "000101010",
                            7230 => "101000000",
                            7231 => "001001110",
                            7232 => "001110110",
                            7233 => "011111010",
                            7234 => "100001110",
                            7235 => "010000000",
                            7236 => "101001100",
                            7237 => "101110010",
                            7238 => "000110100",
                            7239 => "111000010",
                            7240 => "010001110",
                            7241 => "011100010",
                            7242 => "101001010",
                            7243 => "100100000",
                            7244 => "100010100",
                            7245 => "010010110",
                            7246 => "100011100",
                            7247 => "000110000",
                            7248 => "100111000",
                            7249 => "101101100",
                            7250 => "110100000",
                            7251 => "000101110",
                            7252 => "010010110",
                            7253 => "000010010",
                            7254 => "000000000",
                            7255 => "001001110",
                            7256 => "100100000",
                            7257 => "111001100",
                            7258 => "001000010",
                            7259 => "010101110",
                            7260 => "000010000",
                            7261 => "000000000",
                            7262 => "010001011",
                            7263 => "000000000",
                            7264 => "000000000",
                            7265 => "010001000",
                            7266 => "011101110",
                            7267 => "101010100",
                            7268 => "010000000",
                            7269 => "000000000",
                            7270 => "010100010",
                            7271 => "000001100",
                            7272 => "010010100",
                            7273 => "101110000",
                            7274 => "000111110",
                            7275 => "000011010",
                            7276 => "010010000",
                            7277 => "000010000",
                            7278 => "000010100",
                            7279 => "110100010",
                            7280 => "111101010",
                            7281 => "011010110",
                            7282 => "000000010",
                            7283 => "101110110",
                            7284 => "111101000",
                            7285 => "000110110",
                            7286 => "001000010",
                            7287 => "011111010",
                            7288 => "011011100",
                            7289 => "000100100",
                            7290 => "011000010",
                            7291 => "011110100",
                            7292 => "100000010",
                            7293 => "010110110",
                            7294 => "010100000",
                            7295 => "000110000",
                            7296 => "000000010",
                            7297 => "001110100",
                            7298 => "000110000",
                            7299 => "100010010",
                            7300 => "000000000",
                            7301 => "000000000",
                            7302 => "000101110",
                            7303 => "000000110",
                            7304 => "000000110",
                            7305 => "000000000",
                            7306 => "000101110",
                            7307 => "111111010",
                            7308 => "000001000",
                            7309 => "000010110",
                            7310 => "001001010",
                            7311 => "000101010",
                            7312 => "100111110",
                            7313 => "011111110",
                            7314 => "111111110",
                            7315 => "000101110",
                            7316 => "110100100",
                            7317 => "010001000",
                            7318 => "011110110",
                            7319 => "000101000",
                            7320 => "111101110",
                            7321 => "110010010",
                            7322 => "011010010",
                            7323 => "111000110",
                            7324 => "001110100",
                            7325 => "100101100",
                            7326 => "111111000",
                            7327 => "001100010",
                            7328 => "111001100",
                            7329 => "110110000",
                            7330 => "000000000",
                            7331 => "000000000",
                            7332 => "000011000",
                            7333 => "100111110",
                            7334 => "111100100",
                            7335 => "010101110",
                            7336 => "100111000",
                            7337 => "101101100",
                            7338 => "110100000",
                            7339 => "000101110",
                            7340 => "010010110",
                            7341 => "000010010",
                            7342 => "000010000",
                            7343 => "000000000",
                            7344 => "010001011",
                            7345 => "000000000",
                            7346 => "000000000",
                            7347 => "001010000",
                            7348 => "100101010",
                            7349 => "001110100",
                            7350 => "010000000",
                            7351 => "000000000",
                            7352 => "100000000",
                            7353 => "000001100",
                            7354 => "001110010",
                            7355 => "110011110",
                            7356 => "000010100",
                            7357 => "110100010",
                            7358 => "111101010",
                            7359 => "011010110",
                            7360 => "101000100",
                            7361 => "100111110",
                            7362 => "100010000",
                            7363 => "111010100",
                            7364 => "111001110",
                            7365 => "000101110",
                            7366 => "000000010",
                            7367 => "101110110",
                            7368 => "011101110",
                            7369 => "001011010",
                            7370 => "101000110",
                            7371 => "110001100",
                            7372 => "000011110",
                            7373 => "001010110",
                            7374 => "100101100",
                            7375 => "011011110",
                            7376 => "010100000",
                            7377 => "000100000",
                            7378 => "000000010",
                            7379 => "111111010",
                            7380 => "110110000",
                            7381 => "101011110",
                            7382 => "000000000",
                            7383 => "000000000",
                            7384 => "000000000",
                            7385 => "000000000",
                            7386 => "000011000",
                            7387 => "100111110",
                            7388 => "111100100",
                            7389 => "010101110",
                            7390 => "100111000",
                            7391 => "101101100",
                            7392 => "110100000",
                            7393 => "000101110",
                            7394 => "010010110",
                            7395 => "000010010",
                            7396 => "000010000",
                            7397 => "000000000",
                            7398 => "010001011",
                            7399 => "000000000",
                            7400 => "000000000",
                            7401 => "001010000",
                            7402 => "111010000",
                            7403 => "001000110",
                            7404 => "010000000",
                            7405 => "000000000",
                            7406 => "100000000",
                            7407 => "000001100",
                            7408 => "101010110",
                            7409 => "010110100",
                            7410 => "000010100",
                            7411 => "110100010",
                            7412 => "111101010",
                            7413 => "011010110",
                            7414 => "000111110",
                            7415 => "000011010",
                            7416 => "010010000",
                            7417 => "000010000",
                            7418 => "111101000",
                            7419 => "000110110",
                            7420 => "000000010",
                            7421 => "101110110",
                            7422 => "011000010",
                            7423 => "011110100",
                            7424 => "100000010",
                            7425 => "010110110",
                            7426 => "001000010",
                            7427 => "011111010",
                            7428 => "011011100",
                            7429 => "001011100",
                            7430 => "010100000",
                            7431 => "000100000",
                            7432 => "000000010",
                            7433 => "111111000",
                            7434 => "110111100",
                            7435 => "001011100",
                            7436 => "000000000",
                            7437 => "000000000",
                            7438 => "000000000",
                            7439 => "000000000",
                            7440 => "000011000",
                            7441 => "100111110",
                            7442 => "111100100",
                            7443 => "010101110",
                            7444 => "100111000",
                            7445 => "101101100",
                            7446 => "110100000",
                            7447 => "000101110",
                            7448 => "010010110",
                            7449 => "000010010",
                            7450 => "000010000",
                            7451 => "000000000",
                            7452 => "010001011",
                            7453 => "000000000",
                            7454 => "000000000",
                            7455 => "001010000",
                            7456 => "100010100",
                            7457 => "010101110",
                            7458 => "010000000",
                            7459 => "000000000",
                            7460 => "100000000",
                            7461 => "000001100",
                            7462 => "011110000",
                            7463 => "110100010",
                            7464 => "000010100",
                            7465 => "110100010",
                            7466 => "111101010",
                            7467 => "011010110",
                            7468 => "101011000",
                            7469 => "010000110",
                            7470 => "010010110",
                            7471 => "001001110",
                            7472 => "110011000",
                            7473 => "010000010",
                            7474 => "000000010",
                            7475 => "101110110",
                            7476 => "011111010",
                            7477 => "000101000",
                            7478 => "111111110",
                            7479 => "100011000",
                            7480 => "000111110",
                            7481 => "010111110",
                            7482 => "111010000",
                            7483 => "011011010",
                            7484 => "010100000",
                            7485 => "000100010",
                            7486 => "000000010",
                            7487 => "111111100",
                            7488 => "011000110",
                            7489 => "110000110",
                            7490 => "000000000",
                            7491 => "000000000",
                            7492 => "000000000",
                            7493 => "000000000",
                            7494 => "000011000",
                            7495 => "100111110",
                            7496 => "111100100",
                            7497 => "010101110",
                            7498 => "100111000",
                            7499 => "101101100",
                            7500 => "110100000",
                            7501 => "000101110",
                            7502 => "010010110",
                            7503 => "000010010",
                            7504 => "000010000",
                            7505 => "000000000",
                            7506 => "010001011",
                            7507 => "000000000",
                            7508 => "000000000",
                            7509 => "001101000",
                            7510 => "111111010",
                            7511 => "111111110",
                            7512 => "010000000",
                            7513 => "000000000",
                            7514 => "100000000",
                            7515 => "000001100",
                            7516 => "111010000",
                            7517 => "000111110",
                            7518 => "000010100",
                            7519 => "110100010",
                            7520 => "111101010",
                            7521 => "011010110",
                            7522 => "110000000",
                            7523 => "001001100",
                            7524 => "010101000",
                            7525 => "010000010",
                            7526 => "110011000",
                            7527 => "010110100",
                            7528 => "000000000",
                            7529 => "010100000",
                            7530 => "001000110",
                            7531 => "011111100",
                            7532 => "000011010",
                            7533 => "100100010",
                            7534 => "000000000",
                            7535 => "000000000",
                            7536 => "000000000",
                            7537 => "000000000",
                            7538 => "100000000",
                            7539 => "000000100",
                            7540 => "111110100",
                            7541 => "111100000",
                            7542 => "011000010",
                            7543 => "110000010",
                            7544 => "000000000",
                            7545 => "000000000",
                            7546 => "000000100",
                            7547 => "000001000",
                            7548 => "000001010",
                            7549 => "101101000",
                            7550 => "000000010",
                            7551 => "000000110",
                            7552 => "000000110",
                            7553 => "000010000",
                            7554 => "000000010",
                            7555 => "000000010",
                            7556 => "000001000",
                            7557 => "000000100",
                            7558 => "000000000",
                            7559 => "000000000",
                            7560 => "000011000",
                            7561 => "100111110",
                            7562 => "111100100",
                            7563 => "010101110",
                            7564 => "100111000",
                            7565 => "101101100",
                            7566 => "110100000",
                            7567 => "000101110",
                            7568 => "010010110",
                            7569 => "000010010",
                            7570 => "000010000",
                            7571 => "000000000",
                            7572 => "010001011",
                            7573 => "000000000",
                            7574 => "000000000",
                            7575 => "001101000",
                            7576 => "111111100",
                            7577 => "000000000",
                            7578 => "010000000",
                            7579 => "000000000",
                            7580 => "100000000",
                            7581 => "000001100",
                            7582 => "111010000",
                            7583 => "000111100",
                            7584 => "000010100",
                            7585 => "110100010",
                            7586 => "111101010",
                            7587 => "011010110",
                            7588 => "110000000",
                            7589 => "001001100",
                            7590 => "010101000",
                            7591 => "010000010",
                            7592 => "110011000",
                            7593 => "010110110",
                            7594 => "000000000",
                            7595 => "010100000",
                            7596 => "110011110",
                            7597 => "110010110",
                            7598 => "101111100",
                            7599 => "000000110",
                            7600 => "000000000",
                            7601 => "000000000",
                            7602 => "000000000",
                            7603 => "000000000",
                            7604 => "100000000",
                            7605 => "000000100",
                            7606 => "111110100",
                            7607 => "111100000",
                            7608 => "000001010",
                            7609 => "000000000",
                            7610 => "000000000",
                            7611 => "000000000",
                            7612 => "000000100",
                            7613 => "000001000",
                            7614 => "000001010",
                            7615 => "101101000",
                            7616 => "000000010",
                            7617 => "000000110",
                            7618 => "000000110",
                            7619 => "000010000",
                            7620 => "000000010",
                            7621 => "000000010",
                            7622 => "000001000",
                            7623 => "000000100",
                            7624 => "100111000",
                            7625 => "101101100",
                            7626 => "110100000",
                            7627 => "000101110",
                            7628 => "010010110",
                            7629 => "000010010",
                            7630 => "000000000",
                            7631 => "001001110",
                            7632 => "100100000",
                            7633 => "111001100",
                            7634 => "001000010",
                            7635 => "010101110",
                            7636 => "000010000",
                            7637 => "000000000",
                            7638 => "010001011",
                            7639 => "000000000",
                            7640 => "000000000",
                            7641 => "001010000",
                            7642 => "001011000",
                            7643 => "101111010",
                            7644 => "010000000",
                            7645 => "000000000",
                            7646 => "001101000",
                            7647 => "000001100",
                            7648 => "001000100",
                            7649 => "011011000",
                            7650 => "101011000",
                            7651 => "010000110",
                            7652 => "010010110",
                            7653 => "001001110",
                            7654 => "000010100",
                            7655 => "110100010",
                            7656 => "111101010",
                            7657 => "011010110",
                            7658 => "000000010",
                            7659 => "101110110",
                            7660 => "110011000",
                            7661 => "010000010",
                            7662 => "000111110",
                            7663 => "010111110",
                            7664 => "111010000",
                            7665 => "011011010",
                            7666 => "011111010",
                            7667 => "000101000",
                            7668 => "111111110",
                            7669 => "100011010",
                            7670 => "010100000",
                            7671 => "000100010",
                            7672 => "000000000",
                            7673 => "010000100",
                            7674 => "011001010",
                            7675 => "011111100",
                            7676 => "000000000",
                            7677 => "000000000",
                            7678 => "000000000",
                            7679 => "000000000",
                            7680 => "000011000",
                            7681 => "100111110",
                            7682 => "111100100",
                            7683 => "010101110",
                            7684 => "100111000",
                            7685 => "101101100",
                            7686 => "110100000",
                            7687 => "000101110",
                            7688 => "010010110",
                            7689 => "000010010",
                            7690 => "000010000",
                            7691 => "000000000",
                            7692 => "010001011",
                            7693 => "000000000",
                            7694 => "000000000",
                            7695 => "001010000",
                            7696 => "100010100",
                            7697 => "010110000",
                            7698 => "010000000",
                            7699 => "000000000",
                            7700 => "100000000",
                            7701 => "000001100",
                            7702 => "011110000",
                            7703 => "110100000",
                            7704 => "000010100",
                            7705 => "110100010",
                            7706 => "111101010",
                            7707 => "011010110",
                            7708 => "101011000",
                            7709 => "010000110",
                            7710 => "010010110",
                            7711 => "001001110",
                            7712 => "110011000",
                            7713 => "010000010",
                            7714 => "000000010",
                            7715 => "101110110",
                            7716 => "011111010",
                            7717 => "000101000",
                            7718 => "111111110",
                            7719 => "100011010",
                            7720 => "000111110",
                            7721 => "010111110",
                            7722 => "111010000",
                            7723 => "011011100",
                            7724 => "010100000",
                            7725 => "000100000",
                            7726 => "000000010",
                            7727 => "111111100",
                            7728 => "011000110",
                            7729 => "110000100",
                            7730 => "000000000",
                            7731 => "000000000",
                            7732 => "100111000",
                            7733 => "101101100",
                            7734 => "110100000",
                            7735 => "000101110",
                            7736 => "010010110",
                            7737 => "000010010",
                            7738 => "000000000",
                            7739 => "001001110",
                            7740 => "100100000",
                            7741 => "111001100",
                            7742 => "001000010",
                            7743 => "010101110",
                            7744 => "000010000",
                            7745 => "000000000",
                            7746 => "010001011",
                            7747 => "000000000",
                            7748 => "000000000",
                            7749 => "001100000",
                            7750 => "110111110",
                            7751 => "000110110",
                            7752 => "010000000",
                            7753 => "000000000",
                            7754 => "111101110",
                            7755 => "000001100",
                            7756 => "100100000",
                            7757 => "000001110",
                            7758 => "110000000",
                            7759 => "001001100",
                            7760 => "010101000",
                            7761 => "010000010",
                            7762 => "000010100",
                            7763 => "110100010",
                            7764 => "111101010",
                            7765 => "011010110",
                            7766 => "000000000",
                            7767 => "010100000",
                            7768 => "110011000",
                            7769 => "010110110",
                            7770 => "100011000",
                            7771 => "011000000",
                            7772 => "000110000",
                            7773 => "100100010",
                            7774 => "110011110",
                            7775 => "110010110",
                            7776 => "101111100",
                            7777 => "000001000",
                            7778 => "011100000",
                            7779 => "000100100",
                            7780 => "010011100",
                            7781 => "001000000",
                            7782 => "001000100",
                            7783 => "101100000",
                            7784 => "000000000",
                            7785 => "000000000",
                            7786 => "000000100",
                            7787 => "000001000",
                            7788 => "000001000",
                            7789 => "111000100",
                            7790 => "000001000",
                            7791 => "000000100",
                            7792 => "000000000",
                            7793 => "000000000",
                            7794 => "000000000",
                            7795 => "000000000",
                            7796 => "000011000",
                            7797 => "100111110",
                            7798 => "111100100",
                            7799 => "010101110",
                            7800 => "100111000",
                            7801 => "101101100",
                            7802 => "110100000",
                            7803 => "000101110",
                            7804 => "010010110",
                            7805 => "000010010",
                            7806 => "000010000",
                            7807 => "000000000",
                            7808 => "010001011",
                            7809 => "000000000",
                            7810 => "000000000",
                            7811 => "001010000",
                            7812 => "111111100",
                            7813 => "000000010",
                            7814 => "010000000",
                            7815 => "000000000",
                            7816 => "100000000",
                            7817 => "000001100",
                            7818 => "111010000",
                            7819 => "001010010",
                            7820 => "000010100",
                            7821 => "110100010",
                            7822 => "111101010",
                            7823 => "011010110",
                            7824 => "110000000",
                            7825 => "001001100",
                            7826 => "010101000",
                            7827 => "010000010",
                            7828 => "110011000",
                            7829 => "010110110",
                            7830 => "000000000",
                            7831 => "010100000",
                            7832 => "110011110",
                            7833 => "110010110",
                            7834 => "101111100",
                            7835 => "000001000",
                            7836 => "100011000",
                            7837 => "011000000",
                            7838 => "000110000",
                            7839 => "100100100",
                            7840 => "010100000",
                            7841 => "000100000",
                            7842 => "111110100",
                            7843 => "111100000",
                            7844 => "101000000",
                            7845 => "110100000",
                            7846 => "000000000",
                            7847 => "000000000",
                            7848 => "100111000",
                            7849 => "101101100",
                            7850 => "110100000",
                            7851 => "000101110",
                            7852 => "010010110",
                            7853 => "000010010",
                            7854 => "000000000",
                            7855 => "001001110",
                            7856 => "100100000",
                            7857 => "111001100",
                            7858 => "001000010",
                            7859 => "010101110",
                            7860 => "000010000",
                            7861 => "000000000",
                            7862 => "010001011",
                            7863 => "000000000",
                            7864 => "000000000",
                            7865 => "001100000",
                            7866 => "110100100",
                            7867 => "011010000",
                            7868 => "010000000",
                            7869 => "000000000",
                            7870 => "111101110",
                            7871 => "000001100",
                            7872 => "100111000",
                            7873 => "101110100",
                            7874 => "110000000",
                            7875 => "001001100",
                            7876 => "010101000",
                            7877 => "010000010",
                            7878 => "000010100",
                            7879 => "110100010",
                            7880 => "111101010",
                            7881 => "011010110",
                            7882 => "000000000",
                            7883 => "010100000",
                            7884 => "110011000",
                            7885 => "010110100",
                            7886 => "011000100",
                            7887 => "110011100",
                            7888 => "110001100",
                            7889 => "111010110",
                            7890 => "001000110",
                            7891 => "011111100",
                            7892 => "000011010",
                            7893 => "100100100",
                            7894 => "011100000",
                            7895 => "000100100",
                            7896 => "010011100",
                            7897 => "001000000",
                            7898 => "111110100",
                            7899 => "101010000",
                            7900 => "000000000",
                            7901 => "000000000",
                            7902 => "000000100",
                            7903 => "000001000",
                            7904 => "000001000",
                            7905 => "111000100",
                            7906 => "000001000",
                            7907 => "000000100",
                            7908 => "000000000",
                            7909 => "000000000",
                            7910 => "000000000",
                            7911 => "000000000",
                            7912 => "000011000",
                            7913 => "100111110",
                            7914 => "111100100",
                            7915 => "010101110",
                            7916 => "100111000",
                            7917 => "101101100",
                            7918 => "110100000",
                            7919 => "000101110",
                            7920 => "010010110",
                            7921 => "000010010",
                            7922 => "000010000",
                            7923 => "000000000",
                            7924 => "010001011",
                            7925 => "000000000",
                            7926 => "000000000",
                            7927 => "001010000",
                            7928 => "111111100",
                            7929 => "000000100",
                            7930 => "010000000",
                            7931 => "000000000",
                            7932 => "100000000",
                            7933 => "000001100",
                            7934 => "111010000",
                            7935 => "001010000",
                            7936 => "000010100",
                            7937 => "110100010",
                            7938 => "111101010",
                            7939 => "011010110",
                            7940 => "110000000",
                            7941 => "001001100",
                            7942 => "010101000",
                            7943 => "010000010",
                            7944 => "110011000",
                            7945 => "010110100",
                            7946 => "000000000",
                            7947 => "010100000",
                            7948 => "001000110",
                            7949 => "011111100",
                            7950 => "000011010",
                            7951 => "100100100",
                            7952 => "011000100",
                            7953 => "110011100",
                            7954 => "110001100",
                            7955 => "111011000",
                            7956 => "010100000",
                            7957 => "000100000",
                            7958 => "111110100",
                            7959 => "111100000",
                            7960 => "011110000",
                            7961 => "110010010",
                            7962 => "000000000",
                            7963 => "000000000",
                            7964 => "000000000",
                            7965 => "000000000",
                            7966 => "000011000",
                            7967 => "100111110",
                            7968 => "111100100",
                            7969 => "010101110",
                            7970 => "100111000",
                            7971 => "101101100",
                            7972 => "110100000",
                            7973 => "000101110",
                            7974 => "010010110",
                            7975 => "000010010",
                            7976 => "000010000",
                            7977 => "000000000",
                            7978 => "010001011",
                            7979 => "000000000",
                            7980 => "000000110",
                            7981 => "100101100",
                            7982 => "111111100",
                            7983 => "000000110",
                            7984 => "010000000",
                            7985 => "000000000",
                            7986 => "100000000",
                            7987 => "000001100",
                            7988 => "111001000",
                            7989 => "101110010",
                            7990 => "000010100",
                            7991 => "110100010",
                            7992 => "111101010",
                            7993 => "011010110",
                            7994 => "110000000",
                            7995 => "001001100",
                            7996 => "010101000",
                            7997 => "010000010",
                            7998 => "110011000",
                            7999 => "010110110",
                            8000 => "000000000",
                            8001 => "010100000",
                            8002 => "110011110",
                            8003 => "110010110",
                            8004 => "101111100",
                            8005 => "000001000",
                            8006 => "100011000",
                            8007 => "011000000",
                            8008 => "000110000",
                            8009 => "100100100",
                            8010 => "010100000",
                            8011 => "000110000",
                            8012 => "111110100",
                            8013 => "111100000",
                            8014 => "011100010",
                            8015 => "111010110",
                            8016 => "000000000",
                            8017 => "000000000",
                            8018 => "010001110",
                            8019 => "010001010",
                            8020 => "010101000",
                            8021 => "001000000",
                            8022 => "001011110",
                            8023 => "001000000",
                            8024 => "010010000",
                            8025 => "010101000",
                            8026 => "010101000",
                            8027 => "010100000",
                            8028 => "001011110",
                            8029 => "001100010",
                            8030 => "001011100",
                            8031 => "001100010",
                            8032 => "000011010",
                            8033 => "000010100",
                            8034 => "010010000",
                            8035 => "011011110",
                            8036 => "011100110",
                            8037 => "011101000",
                            8038 => "001110100",
                            8039 => "001000000",
                            8040 => "011001000",
                            8041 => "011101000",
                            8042 => "011101010",
                            8043 => "001011100",
                            8044 => "011001000",
                            8045 => "011010110",
                            8046 => "000011010",
                            8047 => "000010100",
                            8048 => "010000110",
                            8049 => "011011110",
                            8050 => "011011100",
                            8051 => "011011100",
                            8052 => "011001010",
                            8053 => "011000110",
                            8054 => "011101000",
                            8055 => "011010010",
                            8056 => "011011110",
                            8057 => "011011100",
                            8058 => "001110100",
                            8059 => "001000000",
                            8060 => "011010110",
                            8061 => "011001010",
                            8062 => "011001010",
                            8063 => "011100000",
                            8064 => "001011010",
                            8065 => "011000010",
                            8066 => "011011000",
                            8067 => "011010010",
                            8068 => "011101100",
                            8069 => "011001010",
                            8070 => "000011010",
                            8071 => "000010100",
                            8072 => "010001000",
                            8073 => "010011100",
                            8074 => "010101000",
                            8075 => "001110100",
                            8076 => "001000000",
                            8077 => "001100010",
                            8078 => "000011010",
                            8079 => "000010100",
                            8080 => "010101010",
                            8081 => "011100000",
                            8082 => "011001110",
                            8083 => "011100100",
                            8084 => "011000010",
                            8085 => "011001000",
                            8086 => "011001010",
                            8087 => "001011010",
                            8088 => "010010010",
                            8089 => "011011100",
                            8090 => "011100110",
                            8091 => "011001010",
                            8092 => "011000110",
                            8093 => "011101010",
                            8094 => "011100100",
                            8095 => "011001010",
                            8096 => "001011010",
                            8097 => "010100100",
                            8098 => "011001010",
                            8099 => "011100010",
                            8100 => "011101010",
                            8101 => "011001010",
                            8102 => "011100110",
                            8103 => "011101000",
                            8104 => "011100110",
                            8105 => "001110100",
                            8106 => "001000000",
                            8107 => "001100010",
                            8108 => "000011010",
                            8109 => "000010100",
                            8110 => "010101010",
                            8111 => "011100110",
                            8112 => "011001010",
                            8113 => "011100100",
                            8114 => "001011010",
                            8115 => "010000010",
                            8116 => "011001110",
                            8117 => "011001010",
                            8118 => "011011100",
                            8119 => "011101000",
                            8120 => "001110100",
                            8121 => "001000000",
                            8122 => "010011010",
                            8123 => "011011110",
                            8124 => "011110100",
                            8125 => "011010010",
                            8126 => "011011000",
                            8127 => "011011000",
                            8128 => "011000010",
                            8129 => "001011110",
                            8130 => "001101010",
                            8131 => "001011100",
                            8132 => "001100000",
                            8133 => "001000000",
                            8134 => "001010000",
                            8135 => "010101110",
                            8136 => "011010010",
                            8137 => "011011100",
                            8138 => "011001000",
                            8139 => "011011110",
                            8140 => "011101110",
                            8141 => "011100110",
                            8142 => "001000000",
                            8143 => "010011100",
                            8144 => "010101000",
                            8145 => "001000000",
                            8146 => "001100010",
                            8147 => "001100000",
                            8148 => "001011100",
                            8149 => "001100000",
                            8150 => "001110110",
                            8151 => "001000000",
                            8152 => "010101110",
                            8153 => "011010010",
                            8154 => "011011100",
                            8155 => "001101100",
                            8156 => "001101000",
                            8157 => "001110110",
                            8158 => "001000000",
                            8159 => "011110000",
                            8160 => "001101100",
                            8161 => "001101000",
                            8162 => "001010010",
                            8163 => "001000000",
                            8164 => "010000010",
                            8165 => "011100000",
                            8166 => "011100000",
                            8167 => "011011000",
                            8168 => "011001010",
                            8169 => "010101110",
                            8170 => "011001010",
                            8171 => "011000100",
                            8172 => "010010110",
                            8173 => "011010010",
                            8174 => "011101000",
                            8175 => "001011110",
                            8176 => "001101010",
                            8177 => "001100110",
                            8178 => "001101110",
                            8179 => "001011100",
                            8180 => "001100110",
                            8181 => "001101100",
                            8182 => "001000000",
                            8183 => "001010000",
                            8184 => "010010110",
                            8185 => "010010000",
                            8186 => "010101000",
                            8187 => "010011010",
                            8188 => "010011000",
                            8189 => "001011000",
                            8190 => "001000000",
                            8191 => "011011000",
                            8192 => "011010010",
                            8193 => "011010110",
                            8194 => "011001010",
                            8195 => "001000000",
                            8196 => "010001110",
                            8197 => "011001010",
                            8198 => "011000110",
                            8199 => "011010110",
                            8200 => "011011110",
                            8201 => "001010010",
                            8202 => "001000000",
                            8203 => "010000110",
                            8204 => "011010000",
                            8205 => "011100100",
                            8206 => "011011110",
                            8207 => "011011010",
                            8208 => "011001010",
                            8209 => "001011110",
                            8210 => "001110010",
                            8211 => "001101010",
                            8212 => "001011100",
                            8213 => "001100000",
                            8214 => "001011100",
                            8215 => "001101000",
                            8216 => "001101100",
                            8217 => "001100110",
                            8218 => "001110000",
                            8219 => "001011100",
                            8220 => "001101010",
                            8221 => "001101000",
                            8222 => "001000000",
                            8223 => "010100110",
                            8224 => "011000010",
                            8225 => "011001100",
                            8226 => "011000010",
                            8227 => "011100100",
                            8228 => "011010010",
                            8229 => "001011110",
                            8230 => "001101010",
                            8231 => "001100110",
                            8232 => "001101110",
                            8233 => "001011100",
                            8234 => "001100110",
                            8235 => "001101100",
                            8236 => "000011010",
                            8237 => "000010100",
                            8238 => "010000010",
                            8239 => "011000110",
                            8240 => "011000110",
                            8241 => "011001010",
                            8242 => "011100000",
                            8243 => "011101000",
                            8244 => "001110100",
                            8245 => "001000000",
                            8246 => "011101000",
                            8247 => "011001010",
                            8248 => "011110000",
                            8249 => "011101000",
                            8250 => "001011110",
                            8251 => "011010000",
                            8252 => "011101000",
                            8253 => "011011010",
                            8254 => "011011000",
                            8255 => "001011000",
                            8256 => "011000010",
                            8257 => "011100000",
                            8258 => "011100000",
                            8259 => "011011000",
                            8260 => "011010010",
                            8261 => "011000110",
                            8262 => "011000010",
                            8263 => "011101000",
                            8264 => "011010010",
                            8265 => "011011110",
                            8266 => "011011100",
                            8267 => "001011110",
                            8268 => "011110000",
                            8269 => "011010000",
                            8270 => "011101000",
                            8271 => "011011010",
                            8272 => "011011000",
                            8273 => "001010110",
                            8274 => "011110000",
                            8275 => "011011010",
                            8276 => "011011000",
                            8277 => "001011000",
                            8278 => "011000010",
                            8279 => "011100000",
                            8280 => "011100000",
                            8281 => "011011000",
                            8282 => "011010010",
                            8283 => "011000110",
                            8284 => "011000010",
                            8285 => "011101000",
                            8286 => "011010010",
                            8287 => "011011110",
                            8288 => "011011100",
                            8289 => "001011110",
                            8290 => "011110000",
                            8291 => "011011010",
                            8292 => "011011000",
                            8293 => "001110110",
                            8294 => "011100010",
                            8295 => "001111010",
                            8296 => "001100000",
                            8297 => "001011100",
                            8298 => "001110010",
                            8299 => "001011000",
                            8300 => "011010010",
                            8301 => "011011010",
                            8302 => "011000010",
                            8303 => "011001110",
                            8304 => "011001010",
                            8305 => "001011110",
                            8306 => "011000010",
                            8307 => "011101100",
                            8308 => "011010010",
                            8309 => "011001100",
                            8310 => "001011000",
                            8311 => "011010010",
                            8312 => "011011010",
                            8313 => "011000010",
                            8314 => "011001110",
                            8315 => "011001010",
                            8316 => "001011110",
                            8317 => "011101110",
                            8318 => "011001010",
                            8319 => "011000100",
                            8320 => "011100000",
                            8321 => "001011000",
                            8322 => "011010010",
                            8323 => "011011010",
                            8324 => "011000010",
                            8325 => "011001110",
                            8326 => "011001010",
                            8327 => "001011110",
                            8328 => "011000010",
                            8329 => "011100000",
                            8330 => "011011100",
                            8331 => "011001110",
                            8332 => "001011000",
                            8333 => "001010100",
                            8334 => "001011110",
                            8335 => "001010100",
                            8336 => "001110110",
                            8337 => "011100010",
                            8338 => "001111010",
                            8339 => "001100000",
                            8340 => "001011100",
                            8341 => "001110000",
                            8342 => "001011000",
                            8343 => "011000010",
                            8344 => "011100000",
                            8345 => "011100000",
                            8346 => "011011000",
                            8347 => "011010010",
                            8348 => "011000110",
                            8349 => "011000010",
                            8350 => "011101000",
                            8351 => "011010010",
                            8352 => "011011110",
                            8353 => "011011100",
                            8354 => "001011110",
                            8355 => "011100110",
                            8356 => "011010010",
                            8357 => "011001110",
                            8358 => "011011100",
                            8359 => "011001010",
                            8360 => "011001000",
                            8361 => "001011010",
                            8362 => "011001010",
                            8363 => "011110000",
                            8364 => "011000110",
                            8365 => "011010000",
                            8366 => "011000010",
                            8367 => "011011100",
                            8368 => "011001110",
                            8369 => "011001010",
                            8370 => "001110110",
                            8371 => "011101100",
                            8372 => "001111010",
                            8373 => "011000100",
                            8374 => "001100110",
                            8375 => "001110110",
                            8376 => "011100010",
                            8377 => "001111010",
                            8378 => "001100000",
                            8379 => "001011100",
                            8380 => "001110010",
                            8381 => "000011010",
                            8382 => "000010100",
                            8383 => "010000010",
                            8384 => "011000110",
                            8385 => "011000110",
                            8386 => "011001010",
                            8387 => "011100000",
                            8388 => "011101000",
                            8389 => "001011010",
                            8390 => "010001010",
                            8391 => "011011100",
                            8392 => "011000110",
                            8393 => "011011110",
                            8394 => "011001000",
                            8395 => "011010010",
                            8396 => "011011100",
                            8397 => "011001110",
                            8398 => "001110100",
                            8399 => "001000000",
                            8400 => "011001110",
                            8401 => "011110100",
                            8402 => "011010010",
                            8403 => "011100000",
                            8404 => "001011000",
                            8405 => "001000000",
                            8406 => "011001000",
                            8407 => "011001010",
                            8408 => "011001100",
                            8409 => "011011000",
                            8410 => "011000010",
                            8411 => "011101000",
                            8412 => "011001010",
                            8413 => "000011010",
                            8414 => "000010100",
                            8415 => "010000010",
                            8416 => "011000110",
                            8417 => "011000110",
                            8418 => "011001010",
                            8419 => "011100000",
                            8420 => "011101000",
                            8421 => "001011010",
                            8422 => "010011000",
                            8423 => "011000010",
                            8424 => "011011100",
                            8425 => "011001110",
                            8426 => "011101010",
                            8427 => "011000010",
                            8428 => "011001110",
                            8429 => "011001010",
                            8430 => "001110100",
                            8431 => "001000000",
                            8432 => "011001010",
                            8433 => "011011100",
                            8434 => "001011010",
                            8435 => "010101010",
                            8436 => "010100110",
                            8437 => "001011000",
                            8438 => "011001010",
                            8439 => "011011100",
                            8440 => "001110110",
                            8441 => "011100010",
                            8442 => "001111010",
                            8443 => "001100000",
                            8444 => "001011100",
                            8445 => "001110010",
                            8446 => "001011000",
                            8447 => "011001000",
                            8448 => "011000010",
                            8449 => "001110110",
                            8450 => "011100010",
                            8451 => "001111010",
                            8452 => "001100000",
                            8453 => "001011100",
                            8454 => "001110000",
                            8455 => "000011010",
                            8456 => "000010100",
                            8457 => "010000110",
                            8458 => "011011110",
                            8459 => "011011110",
                            8460 => "011010110",
                            8461 => "011010010",
                            8462 => "011001010",
                            8463 => "001110100",
                            8464 => "001000000",
                            8465 => "010111110",
                            8466 => "011001110",
                            8467 => "011000010",
                            8468 => "010111110",
                            8469 => "010011010",
                            8470 => "010010100",
                            8471 => "010100110",
                            8472 => "010011100",
                            8473 => "001110000",
                            8474 => "010101110",
                            8475 => "010101110",
                            8476 => "001110010",
                            8477 => "001110010",
                            8478 => "010000100",
                            8479 => "001111010",
                            8480 => "010001110",
                            8481 => "010100110",
                            8482 => "001100010",
                            8483 => "001011100",
                            8484 => "001100010",
                            8485 => "001011100",
                            8486 => "001100010",
                            8487 => "001101100",
                            8488 => "001100110",
                            8489 => "001101010",
                            8490 => "001101100",
                            8491 => "001110000",
                            8492 => "001100010",
                            8493 => "001100010",
                            8494 => "001100110",
                            8495 => "001100000",
                            8496 => "001011100",
                            8497 => "001100010",
                            8498 => "001011100",
                            8499 => "001100010",
                            8500 => "001011100",
                            8501 => "001100010",
                            8502 => "001101100",
                            8503 => "001100110",
                            8504 => "001101010",
                            8505 => "001101100",
                            8506 => "001110000",
                            8507 => "001100010",
                            8508 => "001100010",
                            8509 => "001101010",
                            8510 => "001110010",
                            8511 => "001011100",
                            8512 => "001100000",
                            8513 => "001110110",
                            8514 => "001000000",
                            8515 => "010111110",
                            8516 => "011001110",
                            8517 => "011000010",
                            8518 => "010111110",
                            8519 => "010000110",
                            8520 => "001100110",
                            8521 => "001101000",
                            8522 => "001100010",
                            8523 => "001101100",
                            8524 => "001100010",
                            8525 => "001100010",
                            8526 => "001101000",
                            8527 => "001110000",
                            8528 => "001110000",
                            8529 => "001111010",
                            8530 => "010001110",
                            8531 => "010100110",
                            8532 => "001100010",
                            8533 => "001011100",
                            8534 => "001100010",
                            8535 => "001011100",
                            8536 => "001100010",
                            8537 => "001101100",
                            8538 => "001100110",
                            8539 => "001101100",
                            8540 => "001101110",
                            8541 => "001100010",
                            8542 => "001100010",
                            8543 => "001101010",
                            8544 => "001100110",
                            8545 => "001110010",
                            8546 => "001011100",
                            8547 => "001100010",
                            8548 => "001011100",
                            8549 => "001100000",
                            8550 => "001011100",
                            8551 => "001100010",
                            8552 => "001101100",
                            8553 => "001100110",
                            8554 => "001101100",
                            8555 => "001101110",
                            8556 => "001100010",
                            8557 => "001100010",
                            8558 => "001101010",
                            8559 => "001101000",
                            8560 => "001101000",
                            8561 => "001011100",
                            8562 => "001100000",
                            8563 => "001110110",
                            8564 => "001000000",
                            8565 => "010111110",
                            8566 => "011001110",
                            8567 => "011000010",
                            8568 => "011000110",
                            8569 => "010111110",
                            8570 => "010101010",
                            8571 => "010000010",
                            8572 => "001011010",
                            8573 => "001100010",
                            8574 => "001101000",
                            8575 => "001101100",
                            8576 => "001100000",
                            8577 => "001101000",
                            8578 => "001110010",
                            8579 => "001110010",
                            8580 => "001101000",
                            8581 => "001110000",
                            8582 => "001011010",
                            8583 => "001100010",
                            8584 => "001111010",
                            8585 => "001100010",
                            8586 => "001011100",
                            8587 => "001100010",
                            8588 => "001101100",
                            8589 => "001100110",
                            8590 => "001101100",
                            8591 => "001110010",
                            8592 => "001100000",
                            8593 => "001110000",
                            8594 => "001100000",
                            8595 => "001110000",
                            8596 => "001100000",
                            8597 => "001011100",
                            8598 => "010000110",
                            8599 => "011010100",
                            8600 => "001100000",
                            8601 => "010010110",
                            8602 => "010000110",
                            8603 => "010100010",
                            8604 => "011010010",
                            8605 => "010000010",
                            8606 => "011010000",
                            8607 => "010011010",
                            8608 => "010011110",
                            8609 => "010011010",
                            8610 => "010000100",
                            8611 => "011010000",
                            8612 => "010001000",
                            8613 => "011010000",
                            8614 => "010000010",
                            8615 => "010100100",
                            8616 => "010010010",
                            8617 => "011100110",
                            8618 => "010000010",
                            8619 => "010100000",
                            8620 => "010101100",
                            8621 => "011011010",
                            8622 => "011011000",
                            8623 => "001011010",
                            8624 => "010010000",
                            8625 => "011101010",
                            8626 => "011010010",
                            8627 => "011011100",
                            8628 => "010110100",
                            8629 => "010100100",
                            8630 => "001110010",
                            8631 => "011110100",
                            8632 => "010010000",
                            8633 => "001011010",
                            8634 => "011101010",
                            8635 => "011001010",
                            8636 => "011100110",
                            8637 => "011001010",
                            8638 => "010101110",
                            8639 => "011001110",
                            8640 => "010001010",
                            8641 => "011110010",
                            8642 => "010011110",
                            8643 => "010011110",
                            8644 => "010010100",
                            8645 => "011100010",
                            8646 => "011110010",
                            8647 => "010010000",
                            8648 => "010110100",
                            8649 => "001100010",
                            8650 => "010000100",
                            8651 => "010011110",
                            8652 => "001101100",
                            8653 => "011101010",
                            8654 => "001101000",
                            8655 => "011001100",
                            8656 => "010100100",
                            8657 => "010001110",
                            8658 => "010010100",
                            8659 => "010100100",
                            8660 => "011110010",
                            8661 => "011100000",
                            8662 => "011000110",
                            8663 => "011110010",
                            8664 => "010100110",
                            8665 => "010101000",
                            8666 => "011000100",
                            8667 => "011010100",
                            8668 => "001101000",
                            8669 => "010011000",
                            8670 => "011011100",
                            8671 => "010001010",
                            8672 => "010001000",
                            8673 => "010100010",
                            8674 => "001100010",
                            8675 => "010101110",
                            8676 => "010101010",
                            8677 => "011000010",
                            8678 => "010000010",
                            8679 => "011011110",
                            8680 => "010000110",
                            8681 => "011011110",
                            8682 => "010001010",
                            8683 => "010000010",
                            8684 => "010011000",
                            8685 => "011101110",
                            8686 => "010111110",
                            8687 => "011101110",
                            8688 => "011000110",
                            8689 => "010000100",
                            8690 => "001110110",
                            8691 => "001000000",
                            8692 => "010111110",
                            8693 => "011001110",
                            8694 => "011000010",
                            8695 => "010111110",
                            8696 => "010110000",
                            8697 => "001100000",
                            8698 => "001110010",
                            8699 => "001100000",
                            8700 => "010001010",
                            8701 => "010010100",
                            8702 => "010010000",
                            8703 => "001101100",
                            8704 => "010110100",
                            8705 => "001110010",
                            8706 => "001111010",
                            8707 => "010001110",
                            8708 => "010100110",
                            8709 => "001100010",
                            8710 => "001011100",
                            8711 => "001100010",
                            8712 => "001011100",
                            8713 => "001100010",
                            8714 => "001101100",
                            8715 => "001100110",
                            8716 => "001101110",
                            8717 => "001100000",
                            8718 => "001101100",
                            8719 => "001101010",
                            8720 => "001100110",
                            8721 => "001101000",
                            8722 => "001100000",
                            8723 => "001011100",
                            8724 => "001110010",
                            8725 => "001011100",
                            8726 => "001100010",
                            8727 => "001011100",
                            8728 => "001100010",
                            8729 => "001101100",
                            8730 => "001100110",
                            8731 => "001101110",
                            8732 => "001100000",
                            8733 => "001101100",
                            8734 => "001101110",
                            8735 => "001100100",
                            8736 => "001101100",
                            8737 => "001101110",
                            8738 => "001011100",
                            8739 => "001100000",
                            8740 => "001110110",
                            8741 => "001000000",
                            8742 => "010111110",
                            8743 => "011001110",
                            8744 => "011010010",
                            8745 => "011001000",
                            8746 => "001111010",
                            8747 => "010001110",
                            8748 => "010000010",
                            8749 => "001100010",
                            8750 => "001011100",
                            8751 => "001100100",
                            8752 => "001011100",
                            8753 => "001101000",
                            8754 => "001110010",
                            8755 => "001100010",
                            8756 => "001110010",
                            8757 => "001100000",
                            8758 => "001110000",
                            8759 => "001110010",
                            8760 => "001101100",
                            8761 => "001101110",
                            8762 => "001011100",
                            8763 => "001100010",
                            8764 => "001101100",
                            8765 => "001100110",
                            8766 => "001101110",
                            8767 => "001100100",
                            8768 => "001100110",
                            8769 => "001101110",
                            8770 => "001100100",
                            8771 => "001100100",
                            8772 => "001101100",
                            8773 => "001110110",
                            8774 => "001000000",
                            8775 => "010111110",
                            8776 => "011001110",
                            8777 => "011000010",
                            8778 => "001111010",
                            8779 => "010001110",
                            8780 => "010000010",
                            8781 => "001100010",
                            8782 => "001011100",
                            8783 => "001100010",
                            8784 => "001011100",
                            8785 => "001100010",
                            8786 => "001101000",
                            8787 => "001110000",
                            8788 => "001110000",
                            8789 => "001101000",
                            8790 => "001101010",
                            8791 => "001110000",
                            8792 => "001100110",
                            8793 => "001100000",
                            8794 => "001100010",
                            8795 => "001011100",
                            8796 => "001100010",
                            8797 => "001101100",
                            8798 => "001100110",
                            8799 => "001100010",
                            8800 => "001100000",
                            8801 => "001100000",
                            8802 => "001101100",
                            8803 => "001101110",
                            8804 => "001101110",
                            8805 => "001100100",
                            8806 => "001110110",
                            8807 => "001000000",
                            8808 => "010111110",
                            8809 => "011001110",
                            8810 => "011000110",
                            8811 => "011011000",
                            8812 => "010111110",
                            8813 => "011000010",
                            8814 => "011101010",
                            8815 => "001111010",
                            8816 => "001100010",
                            8817 => "001011100",
                            8818 => "001100010",
                            8819 => "001011100",
                            8820 => "001100010",
                            8821 => "001100110",
                            8822 => "001110000",
                            8823 => "001110000",
                            8824 => "001110000",
                            8825 => "001100100",
                            8826 => "001110010",
                            8827 => "001100100",
                            8828 => "001110000",
                            8829 => "001100100",
                            8830 => "001011100",
                            8831 => "001100010",
                            8832 => "001101100",
                            8833 => "001100110",
                            8834 => "001101110",
                            8835 => "001100100",
                            8836 => "001100110",
                            8837 => "001101110",
                            8838 => "001100100",
                            8839 => "001100100",
                            8840 => "001110000",
                            8841 => "001110110",
                            8842 => "001000000",
                            8843 => "010111110",
                            8844 => "011001110",
                            8845 => "011000010",
                            8846 => "010111110",
                            8847 => "010101000",
                            8848 => "010011100",
                            8849 => "010010000",
                            8850 => "010001100",
                            8851 => "010000110",
                            8852 => "001100100",
                            8853 => "010110010",
                            8854 => "010101110",
                            8855 => "001101000",
                            8856 => "010100010",
                            8857 => "001111010",
                            8858 => "010001110",
                            8859 => "010100110",
                            8860 => "001100010",
                            8861 => "001011100",
                            8862 => "001100010",
                            8863 => "001011100",
                            8864 => "001100010",
                            8865 => "001101100",
                            8866 => "001100110",
                            8867 => "001101110",
                            8868 => "001100100",
                            8869 => "001100110",
                            8870 => "001101110",
                            8871 => "001100100",
                            8872 => "001100100",
                            8873 => "001101010",
                            8874 => "001011100",
                            8875 => "001101010",
                            8876 => "001101000",
                            8877 => "001011100",
                            8878 => "001100010",
                            8879 => "001011100",
                            8880 => "001100010",
                            8881 => "001101100",
                            8882 => "001100110",
                            8883 => "001101110",
                            8884 => "001100100",
                            8885 => "001100110",
                            8886 => "001101110",
                            8887 => "001100100",
                            8888 => "001101000",
                            8889 => "001110000",
                            8890 => "001011100",
                            8891 => "001100000",
                            8892 => "000011010",
                            8893 => "000010100",
                            8894 => "000011010",
                            8895 => "000010100",
                            8896 => "100111000",
                            8897 => "101101100",
                            8898 => "110100000",
                            8899 => "000101110",
                            8900 => "010010110",
                            8901 => "000010010",
                            8902 => "000000000",
                            8903 => "001001110",
                            8904 => "100100000",
                            8905 => "111001100",
                            8906 => "001000010",
                            8907 => "010101110",
                            8908 => "000010000",
                            8909 => "000000000",
                            8910 => "010001011",
                            8911 => "000000000",
                            8912 => "000000000",
                            8913 => "001010000",
                            8914 => "110111110",
                            8915 => "010010110",
                            8916 => "010000000",
                            8917 => "000000000",
                            8918 => "111101110",
                            8919 => "000001100",
                            8920 => "100011110",
                            8921 => "110111110",
                            8922 => "110000000",
                            8923 => "001001100",
                            8924 => "010101000",
                            8925 => "010000010",
                            8926 => "000010100",
                            8927 => "110100010",
                            8928 => "111101010",
                            8929 => "011010110",
                            8930 => "000000000",
                            8931 => "010100000",
                            8932 => "110011000",
                            8933 => "010110110",
                            8934 => "100011000",
                            8935 => "011000000",
                            8936 => "000110000",
                            8937 => "100100100",
                            8938 => "110011110",
                            8939 => "110010110",
                            8940 => "110000010",
                            8941 => "011100100",
                            8942 => "010100000",
                            8943 => "000100000",
                            8944 => "010100010",
                            8945 => "100011100",
                            8946 => "010001100",
                            8947 => "110001010",
                            8948 => "000000000",
                            8949 => "000000000",
                            8950 => "100111000",
                            8951 => "101101100",
                            8952 => "110100000",
                            8953 => "000101110",
                            8954 => "010010110",
                            8955 => "000010010",
                            8956 => "000000000",
                            8957 => "001001110",
                            8958 => "100100000",
                            8959 => "111001100",
                            8960 => "001000010",
                            8961 => "010101110",
                            8962 => "000010000",
                            8963 => "000000000",
                            8964 => "010001011",
                            8965 => "000000000",
                            8966 => "000000100",
                            8967 => "000100010",
                            8968 => "110111110",
                            8969 => "010110100",
                            8970 => "010000000",
                            8971 => "000000000",
                            8972 => "111101110",
                            8973 => "000001100",
                            8974 => "100011010",
                            8975 => "111001110",
                            8976 => "110000000",
                            8977 => "001001100",
                            8978 => "010101000",
                            8979 => "010000010",
                            8980 => "000010100",
                            8981 => "110100010",
                            8982 => "111101010",
                            8983 => "011010110",
                            8984 => "000000000",
                            8985 => "010100000",
                            8986 => "110011000",
                            8987 => "010110110",
                            8988 => "100011000",
                            8989 => "011000000",
                            8990 => "000110000",
                            8991 => "100100100",
                            8992 => "110011110",
                            8993 => "110010110",
                            8994 => "110000010",
                            8995 => "011100100",
                            8996 => "010100000",
                            8997 => "000110000",
                            8998 => "010100010",
                            8999 => "100011100",
                            9000 => "011000100",
                            9001 => "100010010",
                            9002 => "000000000",
                            9003 => "000000000",
                            9004 => "010010000",
                            9005 => "010101000",
                            9006 => "010101000",
                            9007 => "010100000",
                            9008 => "001011110",
                            9009 => "001100010",
                            9010 => "001011100",
                            9011 => "001100010",
                            9012 => "001000000",
                            9013 => "001100110",
                            9014 => "001100000",
                            9015 => "001100100",
                            9016 => "001000000",
                            9017 => "010001100",
                            9018 => "011011110",
                            9019 => "011101010",
                            9020 => "011011100",
                            9021 => "011001000",
                            9022 => "000011010",
                            9023 => "000010100",
                            9024 => "010001000",
                            9025 => "011000010",
                            9026 => "011101000",
                            9027 => "011001010",
                            9028 => "001110100",
                            9029 => "001000000",
                            9030 => "010101000",
                            9031 => "011010000",
                            9032 => "011101010",
                            9033 => "001011000",
                            9034 => "001000000",
                            9035 => "001100010",
                            9036 => "001110000",
                            9037 => "001000000",
                            9038 => "010011100",
                            9039 => "011011110",
                            9040 => "011101100",
                            9041 => "001000000",
                            9042 => "001100100",
                            9043 => "001100000",
                            9044 => "001100100",
                            9045 => "001100010",
                            9046 => "001000000",
                            9047 => "001100010",
                            9048 => "001100100",
                            9049 => "001110100",
                            9050 => "001100100",
                            9051 => "001100010",
                            9052 => "001110100",
                            9053 => "001100000",
                            9054 => "001100000",
                            9055 => "001000000",
                            9056 => "010001110",
                            9057 => "010011010",
                            9058 => "010101000",
                            9059 => "000011010",
                            9060 => "000010100",
                            9061 => "010100110",
                            9062 => "011001010",
                            9063 => "011100100",
                            9064 => "011101100",
                            9065 => "011001010",
                            9066 => "011100100",
                            9067 => "001110100",
                            9068 => "001000000",
                            9069 => "010000010",
                            9070 => "011100000",
                            9071 => "011000010",
                            9072 => "011000110",
                            9073 => "011010000",
                            9074 => "011001010",
                            9075 => "000011010",
                            9076 => "000010100",
                            9077 => "010011000",
                            9078 => "011011110",
                            9079 => "011000110",
                            9080 => "011000010",
                            9081 => "011101000",
                            9082 => "011010010",
                            9083 => "011011110",
                            9084 => "011011100",
                            9085 => "001110100",
                            9086 => "001000000",
                            9087 => "011010000",
                            9088 => "011101000",
                            9089 => "011101000",
                            9090 => "011100000",
                            9091 => "001110100",
                            9092 => "001011110",
                            9093 => "001011110",
                            9094 => "011101110",
                            9095 => "011101110",
                            9096 => "011101110",
                            9097 => "001011100",
                            9098 => "011001000",
                            9099 => "011101000",
                            9100 => "011101010",
                            9101 => "001011100",
                            9102 => "011001000",
                            9103 => "011010110",
                            9104 => "001011110",
                            9105 => "000011010",
                            9106 => "000010100",
                            9107 => "010000110",
                            9108 => "011011110",
                            9109 => "011011100",
                            9110 => "011101000",
                            9111 => "011001010",
                            9112 => "011011100",
                            9113 => "011101000",
                            9114 => "001011010",
                            9115 => "010011000",
                            9116 => "011001010",
                            9117 => "011011100",
                            9118 => "011001110",
                            9119 => "011101000",
                            9120 => "011010000",
                            9121 => "001110100",
                            9122 => "001000000",
                            9123 => "001100100",
                            9124 => "001100000",
                            9125 => "001100100",
                            9126 => "000011010",
                            9127 => "000010100",
                            9128 => "010000110",
                            9129 => "011011110",
                            9130 => "011011100",
                            9131 => "011011100",
                            9132 => "011001010",
                            9133 => "011000110",
                            9134 => "011101000",
                            9135 => "011010010",
                            9136 => "011011110",
                            9137 => "011011100",
                            9138 => "001110100",
                            9139 => "001000000",
                            9140 => "011000110",
                            9141 => "011011000",
                            9142 => "011011110",
                            9143 => "011100110",
                            9144 => "011001010",
                            9145 => "000011010",
                            9146 => "000010100",
                            9147 => "010000110",
                            9148 => "011011110",
                            9149 => "011011100",
                            9150 => "011101000",
                            9151 => "011001010",
                            9152 => "011011100",
                            9153 => "011101000",
                            9154 => "001011010",
                            9155 => "010101000",
                            9156 => "011110010",
                            9157 => "011100000",
                            9158 => "011001010",
                            9159 => "001110100",
                            9160 => "001000000",
                            9161 => "011101000",
                            9162 => "011001010",
                            9163 => "011110000",
                            9164 => "011101000",
                            9165 => "001011110",
                            9166 => "011010000",
                            9167 => "011101000",
                            9168 => "011011010",
                            9169 => "011011000",
                            9170 => "001110110",
                            9171 => "001000000",
                            9172 => "011000110",
                            9173 => "011010000",
                            9174 => "011000010",
                            9175 => "011100100",
                            9176 => "011100110",
                            9177 => "011001010",
                            9178 => "011101000",
                            9179 => "001111010",
                            9180 => "011010010",
                            9181 => "011100110",
                            9182 => "011011110",
                            9183 => "001011010",
                            9184 => "001110000",
                            9185 => "001110000",
                            9186 => "001101010",
                            9187 => "001110010",
                            9188 => "001011010",
                            9189 => "001100010",
                            9190 => "000011010",
                            9191 => "000010100",
                            9192 => "010100110",
                            9193 => "011001010",
                            9194 => "011101000",
                            9195 => "001011010",
                            9196 => "010000110",
                            9197 => "011011110",
                            9198 => "011011110",
                            9199 => "011010110",
                            9200 => "011010010",
                            9201 => "011001010",
                            9202 => "001110100",
                            9203 => "001000000",
                            9204 => "010000100",
                            9205 => "010010010",
                            9206 => "010001110",
                            9207 => "011010010",
                            9208 => "011100000",
                            9209 => "010100110",
                            9210 => "011001010",
                            9211 => "011100100",
                            9212 => "011101100",
                            9213 => "011001010",
                            9214 => "011100100",
                            9215 => "011111100",
                            9216 => "010000100",
                            9217 => "010010010",
                            9218 => "010101000",
                            9219 => "001011010",
                            9220 => "010010010",
                            9221 => "010100110",
                            9222 => "010001110",
                            9223 => "011111100",
                            9224 => "011100000",
                            9225 => "011011110",
                            9226 => "011011110",
                            9227 => "011011000",
                            9228 => "001011010",
                            9229 => "011100100",
                            9230 => "011001010",
                            9231 => "011001000",
                            9232 => "011010010",
                            9233 => "011100100",
                            9234 => "011001010",
                            9235 => "011000110",
                            9236 => "011101000",
                            9237 => "001011100",
                            9238 => "011000010",
                            9239 => "011010010",
                            9240 => "011101000",
                            9241 => "001011100",
                            9242 => "011001000",
                            9243 => "011101000",
                            9244 => "011101010",
                            9245 => "001011100",
                            9246 => "011001000",
                            9247 => "011010110",
                            9248 => "001111010",
                            9249 => "001101000",
                            9250 => "001100100",
                            9251 => "001101010",
                            9252 => "001101000",
                            9253 => "001100000",
                            9254 => "001101000",
                            9255 => "001100000",
                            9256 => "001110010",
                            9257 => "001101100",
                            9258 => "001011100",
                            9259 => "001100100",
                            9260 => "001100000",
                            9261 => "001101000",
                            9262 => "001110000",
                            9263 => "001100000",
                            9264 => "001011100",
                            9265 => "001100000",
                            9266 => "001100000",
                            9267 => "001100000",
                            9268 => "001100000",
                            9269 => "001110110",
                            9270 => "001000000",
                            9271 => "011100000",
                            9272 => "011000010",
                            9273 => "011101000",
                            9274 => "011010000",
                            9275 => "001111010",
                            9276 => "001011110",
                            9277 => "001110110",
                            9278 => "001000000",
                            9279 => "010010000",
                            9280 => "011101000",
                            9281 => "011101000",
                            9282 => "011100000",
                            9283 => "011011110",
                            9284 => "011011100",
                            9285 => "011011000",
                            9286 => "011110010",
                            9287 => "000011010",
                            9288 => "000010100",
                            9289 => "000011010",
                            9290 => "000010100",
                            9291 => "001111000",
                            9292 => "001000010",
                            9293 => "010001000",
                            9294 => "010011110",
                            9295 => "010000110",
                            9296 => "010101000",
                            9297 => "010110010",
                            9298 => "010100000",
                            9299 => "010001010",
                            9300 => "001000000",
                            9301 => "010010000",
                            9302 => "010101000",
                            9303 => "010011010",
                            9304 => "010011000",
                            9305 => "001000000",
                            9306 => "010100000",
                            9307 => "010101010",
                            9308 => "010000100",
                            9309 => "010011000",
                            9310 => "010010010",
                            9311 => "010000110",
                            9312 => "001000000",
                            9313 => "001000100",
                            9314 => "001011010",
                            9315 => "001011110",
                            9316 => "001011110",
                            9317 => "010010010",
                            9318 => "010001010",
                            9319 => "010101000",
                            9320 => "010001100",
                            9321 => "001011110",
                            9322 => "001011110",
                            9323 => "010001000",
                            9324 => "010101000",
                            9325 => "010001000",
                            9326 => "001000000",
                            9327 => "010010000",
                            9328 => "010101000",
                            9329 => "010011010",
                            9330 => "010011000",
                            9331 => "001000000",
                            9332 => "001100100",
                            9333 => "001011100",
                            9334 => "001100000",
                            9335 => "001011110",
                            9336 => "001011110",
                            9337 => "010001010",
                            9338 => "010011100",
                            9339 => "001000100",
                            9340 => "001111100",
                            9341 => "000010100",
                            9342 => "001111000",
                            9343 => "011010000",
                            9344 => "011101000",
                            9345 => "011011010",
                            9346 => "011011000",
                            9347 => "001111100",
                            9348 => "001111000",
                            9349 => "011010000",
                            9350 => "011001010",
                            9351 => "011000010",
                            9352 => "011001000",
                            9353 => "001111100",
                            9354 => "000010100",
                            9355 => "001111000",
                            9356 => "011101000",
                            9357 => "011010010",
                            9358 => "011101000",
                            9359 => "011011000",
                            9360 => "011001010",
                            9361 => "001111100",
                            9362 => "001100110",
                            9363 => "001100000",
                            9364 => "001100100",
                            9365 => "001000000",
                            9366 => "010001100",
                            9367 => "011011110",
                            9368 => "011101010",
                            9369 => "011011100",
                            9370 => "011001000",
                            9371 => "001111000",
                            9372 => "001011110",
                            9373 => "011101000",
                            9374 => "011010010",
                            9375 => "011101000",
                            9376 => "011011000",
                            9377 => "011001010",
                            9378 => "001111100",
                            9379 => "000010100",
                            9380 => "001111000",
                            9381 => "001011110",
                            9382 => "011010000",
                            9383 => "011001010",
                            9384 => "011000010",
                            9385 => "011001000",
                            9386 => "001111100",
                            9387 => "001111000",
                            9388 => "011000100",
                            9389 => "011011110",
                            9390 => "011001000",
                            9391 => "011110010",
                            9392 => "001111100",
                            9393 => "000010100",
                            9394 => "001111000",
                            9395 => "011010000",
                            9396 => "001100010",
                            9397 => "001111100",
                            9398 => "010001100",
                            9399 => "011011110",
                            9400 => "011101010",
                            9401 => "011011100",
                            9402 => "011001000",
                            9403 => "001111000",
                            9404 => "001011110",
                            9405 => "011010000",
                            9406 => "001100010",
                            9407 => "001111100",
                            9408 => "000010100",
                            9409 => "001111000",
                            9410 => "011100000",
                            9411 => "001111100",
                            9412 => "010101000",
                            9413 => "011010000",
                            9414 => "011001010",
                            9415 => "001000000",
                            9416 => "011001000",
                            9417 => "011011110",
                            9418 => "011000110",
                            9419 => "011101010",
                            9420 => "011011010",
                            9421 => "011001010",
                            9422 => "011011100",
                            9423 => "011101000",
                            9424 => "001000000",
                            9425 => "011010000",
                            9426 => "011000010",
                            9427 => "011100110",
                            9428 => "001000000",
                            9429 => "011011010",
                            9430 => "011011110",
                            9431 => "011101100",
                            9432 => "011001010",
                            9433 => "011001000",
                            9434 => "001000000",
                            9435 => "001111000",
                            9436 => "011000010",
                            9437 => "001000000",
                            9438 => "011010000",
                            9439 => "011100100",
                            9440 => "011001010",
                            9441 => "011001100",
                            9442 => "001111010",
                            9443 => "001000100",
                            9444 => "011010000",
                            9445 => "011101000",
                            9446 => "011101000",
                            9447 => "011100000",
                            9448 => "001110100",
                            9449 => "001011110",
                            9450 => "001011110",
                            9451 => "011101110",
                            9452 => "011101110",
                            9453 => "011101110",
                            9454 => "001011100",
                            9455 => "011001000",
                            9456 => "011101000",
                            9457 => "011101010",
                            9458 => "001011100",
                            9459 => "011001000",
                            9460 => "011010110",
                            9461 => "001011110",
                            9462 => "001000100",
                            9463 => "001111100",
                            9464 => "011010000",
                            9465 => "011001010",
                            9466 => "011100100",
                            9467 => "011001010",
                            9468 => "001111000",
                            9469 => "001011110",
                            9470 => "011000010",
                            9471 => "001111100",
                            9472 => "001011100",
                            9473 => "001111000",
                            9474 => "001011110",
                            9475 => "011100000",
                            9476 => "001111100",
                            9477 => "000010100",
                            9478 => "001111000",
                            9479 => "001011110",
                            9480 => "011000100",
                            9481 => "011011110",
                            9482 => "011001000",
                            9483 => "011110010",
                            9484 => "001111100",
                            9485 => "001111000",
                            9486 => "001011110",
                            9487 => "011010000",
                            9488 => "011101000",
                            9489 => "011011010",
                            9490 => "011011000",
                            9491 => "001111100",
                            9492 => "100111000",
                            9493 => "101101100",
                            9494 => "110100000",
                            9495 => "000101110",
                            9496 => "010010110",
                            9497 => "000010010",
                            9498 => "000000000",
                            9499 => "001001110",
                            9500 => "100100000",
                            9501 => "111001100",
                            9502 => "001000010",
                            9503 => "010101110",
                            9504 => "000010000",
                            9505 => "000000000",
                            9506 => "010001011",
                            9507 => "000000000",
                            9508 => "000000000",
                            9509 => "001010000",
                            9510 => "110111110",
                            9511 => "010111010",
                            9512 => "010000000",
                            9513 => "000000000",
                            9514 => "111101110",
                            9515 => "000001100",
                            9516 => "100011110",
                            9517 => "110011010",
                            9518 => "110000000",
                            9519 => "001001100",
                            9520 => "010101000",
                            9521 => "010000010",
                            9522 => "000010100",
                            9523 => "110100010",
                            9524 => "111101010",
                            9525 => "011010110",
                            9526 => "000000000",
                            9527 => "010100000",
                            9528 => "110011000",
                            9529 => "010110110",
                            9530 => "100011000",
                            9531 => "011000000",
                            9532 => "000110100",
                            9533 => "011110110",
                            9534 => "110011110",
                            9535 => "110010110",
                            9536 => "110000010",
                            9537 => "011100100",
                            9538 => "010100000",
                            9539 => "000100010",
                            9540 => "010100010",
                            9541 => "100011100",
                            9542 => "010001000",
                            9543 => "110110110",
                            9544 => "000000000",
                            9545 => "000000000",
                            9546 => "000000000",
                            9547 => "000000000",
                            9548 => "000011000",
                            9549 => "100111110",
                            9550 => "111100100",
                            9551 => "010101110",
                            9552 => "100111000",
                            9553 => "101101100",
                            9554 => "110100000",
                            9555 => "000101110",
                            9556 => "010010110",
                            9557 => "000010010",
                            9558 => "000010000",
                            9559 => "000000000",
                            9560 => "010001011",
                            9561 => "000000000",
                            9562 => "000000000",
                            9563 => "001010000",
                            9564 => "111111100",
                            9565 => "000001000",
                            9566 => "010000000",
                            9567 => "000000000",
                            9568 => "100000000",
                            9569 => "000001100",
                            9570 => "111010000",
                            9571 => "001001100",
                            9572 => "000010100",
                            9573 => "110100010",
                            9574 => "111101010",
                            9575 => "011010110",
                            9576 => "110000000",
                            9577 => "001001100",
                            9578 => "010101000",
                            9579 => "010000010",
                            9580 => "110011000",
                            9581 => "010110110",
                            9582 => "000000000",
                            9583 => "010100000",
                            9584 => "110011110",
                            9585 => "110010110",
                            9586 => "110000010",
                            9587 => "011100100",
                            9588 => "100011000",
                            9589 => "011000000",
                            9590 => "000110000",
                            9591 => "100100100",
                            9592 => "010100000",
                            9593 => "000100000",
                            9594 => "111110100",
                            9595 => "111100000",
                            9596 => "100111010",
                            9597 => "011000100",
                            9598 => "000000000",
                            9599 => "000000000",
                            9600 => "000000000",
                            9601 => "000000000",
                            9602 => "000011000",
                            9603 => "100111110",
                            9604 => "111100100",
                            9605 => "010101110",
                            9606 => "100111000",
                            9607 => "101101100",
                            9608 => "110100000",
                            9609 => "000101110",
                            9610 => "010010110",
                            9611 => "000010010",
                            9612 => "000010000",
                            9613 => "000000000",
                            9614 => "010001011",
                            9615 => "000000000",
                            9616 => "000000000",
                            9617 => "001010000",
                            9618 => "111111100",
                            9619 => "000001010",
                            9620 => "010000000",
                            9621 => "000000000",
                            9622 => "100000000",
                            9623 => "000001100",
                            9624 => "111010000",
                            9625 => "001001010",
                            9626 => "000010100",
                            9627 => "110100010",
                            9628 => "111101010",
                            9629 => "011010110",
                            9630 => "110000000",
                            9631 => "001001100",
                            9632 => "010101000",
                            9633 => "010000010",
                            9634 => "110011000",
                            9635 => "010110110",
                            9636 => "000000000",
                            9637 => "010100000",
                            9638 => "110011110",
                            9639 => "110010110",
                            9640 => "110000010",
                            9641 => "011100100",
                            9642 => "100011000",
                            9643 => "011000000",
                            9644 => "000110100",
                            9645 => "011111000",
                            9646 => "010100000",
                            9647 => "000100000",
                            9648 => "111110010",
                            9649 => "000001110",
                            9650 => "100111010",
                            9651 => "011000010",
                            9652 => "000000000",
                            9653 => "000000000",
                            9654 => "000000000",
                            9655 => "000000000",
                            9656 => "000011000",
                            9657 => "100111110",
                            9658 => "111100100",
                            9659 => "010101110",
                            9660 => "100111000",
                            9661 => "101101100",
                            9662 => "110100000",
                            9663 => "000101110",
                            9664 => "010010110",
                            9665 => "000010010",
                            9666 => "000010000",
                            9667 => "000000000",
                            9668 => "010001011",
                            9669 => "000000000",
                            9670 => "000000000",
                            9671 => "001010000",
                            9672 => "111111100",
                            9673 => "000001100",
                            9674 => "010000000",
                            9675 => "000000000",
                            9676 => "100000000",
                            9677 => "000001100",
                            9678 => "111010000",
                            9679 => "001001000",
                            9680 => "000010100",
                            9681 => "110100010",
                            9682 => "111101010",
                            9683 => "011010110",
                            9684 => "110000000",
                            9685 => "001001100",
                            9686 => "010101000",
                            9687 => "010000010",
                            9688 => "110011000",
                            9689 => "010110110",
                            9690 => "000000000",
                            9691 => "010100000",
                            9692 => "110011110",
                            9693 => "110010110",
                            9694 => "110000010",
                            9695 => "011100100",
                            9696 => "100011000",
                            9697 => "011000000",
                            9698 => "000110100",
                            9699 => "011111000",
                            9700 => "010100000",
                            9701 => "000100010",
                            9702 => "111110010",
                            9703 => "000001110",
                            9704 => "100111010",
                            9705 => "011000000",
                            9706 => "000000000",
                            9707 => "000000000");

BEGIN
  data_out <= ROM(to_integer(unsigned(address)));
END ARCHITECTURE;

