library IEEE;
library std;
use IEEE.std_logic_1164.all;
use IEEE.NUMERIC_STD.all;

entity delete_keys_rom is
  port (
    address : in std_logic_vector(15 downto 0);
    data_out : out std_logic_vector(8 downto 0) 
  );
end entity;


architecture delete_keys_rom_arch of delete_keys_rom is
type ROM_type is array (0 to 4) of std_logic_vector(95 downto 0);

constant ROM : ROM_type := (
   0 => "111111010110001000101110110000001010100000000001011001100000000110111011111001001111000010111100",
   1 => "111100110001100101000110110000001010100000000001011001100000000110111011111001001110111100100100",
   2 => "110011001111010001110101110000001010100000000001011001100000000110111011111001001111000100001001",
   3 => "000100001001010001000000110000001010100000000001011001100000000110111011111001010000100110010001",
   4 => "001000011000101100001101110000001010100000000001011001100000000110111011111001010001100111001010");

   begin
    data_out <= ROM(to_integer(unsigned(unsigned(address))));
  end architecture;