library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use ieee.math_real.all;

entity Cuckoo_Hashing_tb is
end Cuckoo_Hashing_tb ;

architecture Cuckoo_Hashing_arch of Cuckoo_Hashing_tb is



begin



end architecture ; -- Cuckoo_Hashing_arch
