library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use ieee.math_real.all;

entity SRAM is
  port (
    clock
  ) ;
end SRAM ;

architecture SRAM_arch of SRAM is



begin



end architecture ; -- SRAM_arch
