entity test is

end entity;