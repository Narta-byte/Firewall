library IEEE;
library std;
use IEEE.std_logic_1164.all;
use IEEE.NUMERIC_STD.all;

entity prog_keys_rom is
  port (
    address : in std_logic_vector(6 downto 0);
    data_out : out std_logic_vector(95 downto 0) 
  );
end entity;


architecture prog_keys_rom_arch of prog_keys_rom is
type ROM_type is array (0 to 86) of std_logic_vector(95 downto 0);

constant ROM : ROM_type := (
   0 => "111011010110111011000111110000001010100000000001011001100000000110111011111001001100010110111111",
   1 => "111011010110111011000111110000001010100000000001011001100000000110111011111001001100011011101101",
   2 => "011010111111011000101100110000001010100000000001011001100000000110111011111001001100011100111011",
   3 => "100111110101000010000000110000001010100000000001011001100001111110011100111001001100100010101000",
   4 => "110001101010111011000000110000001010100000000001011001100000000110111011111001001100100111001111",
   5 => "110001101010111011010000110000001010100000000001011001100000000110111011111001001100101001111010",
   6 => "100111110101000010000000110000001010100000000001011001100001111110011100111001001100101110001101",
   7 => "111110110000100110011101110000001010100000000001011001100000000110111011111001001100110111010110",
   8 => "110110000110110101101011110000001010100000000001011001100000000110111011111001001100110011101000",
   9 => "000100101011101000111001110000001010100000000001011001100000000110111011111001001100111011010110",
   10 => "100111110101000010000000110000001010100000000001011001100001111110011100111001001100111111100110",
   11 => "110011001111010001111001110000001010100000000001011001100000000110111011111001001101001100001011",
   12 => "000100001010111100001010110000001010100000000001011001100000000110111011111001001101001010101100",
   13 => "110011001111010000001010110000001010100000000001011001100000000110111011111001001101010001101000",
   14 => "110011001111010000001010110000001010100000000001011001100000000110111011111001001101010001101000",
   15 => "010001111011011100011100110000001010100000000001011001100000000110111011111001001101000001010101",
   16 => "010001111011011100011100110000001010100000000001011001100000000110111011111001001101000100001011",
   17 => "110110010001001101000010110000001010100000000001011001100000000110111011111001001101010110001100",
   18 => "101010110011010100101001110000001010100000000001011001100000000110111011111001001101011000011101",
   19 => "101001011001101111110010110000001010100000000001011001100000000110111011111001001101011110110101",
   20 => "101011000111101001110100110000001010100000000001011001100000000110111011111001001101100011100000",
   21 => "100111110101000010000000110000001010100000000001011001100001111110011100111001001101100111000001",
   22 => "011010110001010111001000110000001010100000000001011001100000000110111011111001001101101010010110",
   23 => "011110011110110100101001110000001010100000000001011001100000000110111011111001001101101100100101",
   24 => "000101101110111000001001110000001010100000000001011001100000000110111011111001001101110001001001",
   25 => "000101101110111000001001110000001010100000000001011001100000000110111011111001001101111011010001",
   26 => "101011000111101001110100110000001010100000000001011001100000000110111011111001001101110101111110",
   27 => "001000010010001110111100110000001010100000000001011001100000000110111011111001001101111111111101",
   28 => "000000000100110100101000110000001010100000000001011001100000000110111011111001001110000010011011",
   29 => "001000011001100001001000110000001010100000000001011001100000000110111011111001001110000101001010",
   30 => "010110100100010100001000110000001010100000000001011001100000000110111011111001001110001001011100",
   31 => "110010010011001001100101110000001010100000000001011001100000000110111011111001001110010101111001",
   32 => "101111000101111111100101110000001010100000000001011001100000000110111011111001001110011011000011",
   33 => "110011001111010000001010110000001010100000000001011001100000000110111011111001001110011100110100",
   34 => "011010110010101000001110110000001010100000000001011001100000000110111011111001001110100010001111",
   35 => "111101001010111001000100110000001010100000000001011001100000000110111011111001001110101010001001",
   36 => "111001010000001001100101110000001010100000000001011001100000000110111011111001001110100100010110",
   37 => "100011100111001000000010110000001010100000000001011001100000000110111011111001001110110010000100",
   38 => "000100010110100101111011110000001010100000000001011001100000000110111011111001001110110100000100",
   39 => "010011001010111001000010110000001010100000000001011001100000000110111011111001001110101100010111",
   40 => "111010000010101011011001110000001010100000000001011001100000000110111011111001001110111010011011",
   41 => "111111010110001000101110110000001010100000000001011001100000000110111011111001001111000010111100",
   42 => "111100110001100101000110110000001010100000000001011001100000000110111011111001001110111100100100",
   43 => "110011001111010001110101110000001010100000000001011001100000000110111011111001001111000100001001",
   44 => "001000011001100001011100110000001010100000000001011001100000000110111011111001001111001000001110",
   45 => "100010111000000000001011110000001010100000000001011001100000000110111011111001001111001100001011",
   46 => "111111010110001000110000110000001010100000000001011001100000000110111011111001001111010010010100",
   47 => "111111010110001000101110110000001010100000000001011001100000000110111011111001001111010100010101",
   48 => "111100010110110101111010110000001010100000000001011001100000000110111011111001001111011010100001",
   49 => "111010000010101011011001110000001010100000000001011001100000000110111011111001001111011100001001",
   50 => "111001011111000001001110110000001010100000000001011001100000000110111011111001001111100010000000",
   51 => "111010000010101000110001110000001010100000000001011001100000000110111011111001001111100100001100",
   52 => "000110100000111010001110110000001010100000000001011001100000000110111011111001001111101011110100",
   53 => "110011001111010001001100110000001010100000000001011001100000000110111011111001001111101100001010",
   54 => "101111000101111111100101110000001010100000000001011001100000000110111011111001001111110000001111",
   55 => "110001110110111010011010110000001010100000000001011001100000000110111011111001001111110111001011",
   56 => "010100100111100100000011110000001010100000000001011001100000000110111011111001001111111010000001",
   57 => "100111001101101000000111110000001010100000000001011001100000000110111011111001001111111111011100",
   58 => "000000001010000000010001110000001010100000000001011001100000000110111011111001010000000010100000",
   59 => "000000001010000000010001110000001010100000000001011001100000000110111011111001010000000101111001",
   60 => "001100110101100010011110110000001010100000000001011001100000000110111011111001010000001010001101",
   61 => "111000000101011000000000110000001010100000000001011001100000000110111011111001010000010000000001",
   62 => "000100101100000111000010110000001010100000000001011001100000000110111011111001010000001100110100",
   63 => "001000011001100000110110110000001010100000000001011001100000000110111011111001010000010110101011",
   64 => "010111100001101100010110110000001010100000000001011001100000000110111011111001010000011001100100",
   65 => "110001110110111010011010110000001010100000000001011001100000000110111011111001010000011101001111",
   66 => "110001110110110010000101110000001010100000000001011001100000000110111011111001010000100000101011",
   67 => "000100001001010001000000110000001010100000000001011001100000000110111011111001010000100110010001",
   68 => "000100001001010001000000110000001010100000000001011001100000000110111011111001010000101001010101",
   69 => "001000011001100001110100110000001010100000000001011001100000000110111011111001010000101100010010",
   70 => "110011001111010001001101110000001010100000000001011001100000000110111011111001010000110011111000",
   71 => "110011001111010001001101110000001010100000000001011001100000000110111011111001010000110011111000",
   72 => "010100011010111111001100110000001010100000000001011001100000000110111011111001010000110110101111",
   73 => "001000000010000111010100110000001010100000000001011001100000000110111011111001010000111001111011",
   74 => "001000000010000111010100110000001010100000000001011001100000000110111011111001010000111110111001",
   75 => "001000011001100001110101110000001010100000000001011001100000000110111011111001010001000010100000",
   76 => "001000011001100001110101110000001010100000000001011001100000000110111011111001010001000010100000",
   77 => "001001100101010000100101110000001010100000000001011001100000000110111011111001010001000111110001",
   78 => "010100100111001000011010110000001010100000000001011001100000000110111011111001010001001000010100",
   79 => "001001100101010000100101110000001010100000000001011001100000000110111011111001010001001111010111",
   80 => "111010000010101011011001110000001010100000000001011001100000000110111011111001010001010001101011",
   81 => "010100100111100100000101110000001010100000000001011001100000000110111011111001010001010111111001",
   82 => "001001100101010000100101110000001010100000000001011001100000000110111011111001010001011011010000",
   83 => "000110100000010011001100110000001010100000000001011001100000000110111011111001010001011101010110",
   84 => "001000011001100001110101110000001010100000000001011001100000000110111011111001010001100011111111",
   85 => "001000011000101100001101110000001010100000000001011001100000000110111011111001010001100111001010",
   86 => "000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000");

   begin
    data_out <= ROM(to_integer(unsigned(unsigned(address))));
  end architecture;


